BZh91AY&SY�؈.��_�ryg����������b�8���T���%J�
�
IUR���J(U)B�*T�URkT�z�I�  
����U%DHT� � I>��  
 P   ( 
(  �y!*�%%  �R$*�B�		)@�UQ$� �pdTP�J�%
��B���
Q��A@a�
� ��!(H��H �(U(� ��   ��
R�� ����� H ��6� �� q@� 	 m�M� -c@:	T)*W�eT�6%UP�L���`y캕UI15�����*I�㪅@�5R
04�u*��bjJ��e��5
(���	R0  @�P�X   ��� ���Vƪ���
�U3j)n�u"��u�QV	[�������(�Q+u�T�ʕq1R(��g+�-�� �wp��9EP����m
����8�`P-�Ҁ� � � n� 6l��k� d � �   m	QX P �)Nz� H �` H   �l
v n��@ ��t8�2H:� ۸QJ
(���46��-� ���A�X ��f@@ � @ � �  1�	�  �Rs� �F�6�4	� G��4� v �
� ��`���ӻ vU$�!
��
4 @��h�X  ��\ A���� ;�4 SF    i$�   �"^yx 9 #�� ` ���� � M�op �`�6� H�@��@�x��{: � ;`l� � ف�d���l��� � " �" ����,ʴ�&�                                    kY�ӈ�������I�       ��������#	���i��4��a"B4?#F��=I�dh���$�(���A�0���&A�F� �� L�S@�*���OI悙4�F � ��D�="���<��� 5 a�F����������'��W��X�͆C<]D��_/�_f���DQ\���(?�AEx�@hE0� ���UE���,|��I]UB:���[4�ϧ���t����g�����|��mG�L���ty�d8��~zq��DXJ��pW�ɉ����|Mc��ʹδ:o�����)�<��lln�Ͷ�x-���l�>��o������� Qt0G�TDA�(v/������ym�3���^\8���zs���oV�e}�bA�[m�Y�
-��(U|�@��g�1�t�iqq��{����/���s-_*�H~/9B
TT�I�
G�,���m�;�S]c��m1��ðI|E_*���B*�U|¿���	���P�R��$�P�_+��A���{ٞqǎ�ƚx�/��i���zy����lS���<Sŗǽ�G��7��4��i�����2��_Ed�+_Ih�搡!R���G�����<Y��n61��{N�8�_T�k����f&@,A�_5i��$�2��5��?�"��AT6��7�>�:{��'���6�����O{��إ��/�_{�|x��)eK�a�[�ھM|�	/�A�_� �z{c�Om6�=q������R��=��g���q�`�c�����}�}�	�B��W��bC_;�ϯc8���m��3�����{����[vI/�����A��?T��,�����F�1�� �|���A������7����Ɖ�َ��;�R���ocot�]u���P�CB�)��շ���$_ C���}q}���m�loi��Ə��m�Pv�o��]���HT��|�LTiZب/��Э��*B���iw����㽦)}���OǶ5�i�`(A¾�ȾQ|���mvP�T6����j /��,�*�H[>��+�@s,b�������HT��Xƾ����h�|���Zx��w��}q�e��&����m����*{�mqOi�S�b�XiB����b$o�ҰX ��B�`��Ǽ�e,�)�<2�v��lm���Ln�x���ciJ{i�@���/�j
���|�`��㽧�M,�O{�=�鱷��)�g��$-��h6�%�Z�bK��U��/� �m��m��a�9rL��|h_/�Pa/������*�U}(B���Ta�l�Z��}�{N�oc�R�Oy�����hP�����A$��c���|�Ɖ޽/{��6���R��7�n/��x���'oM���w������ocm��)J��_i��+���� @��H$�N����ms������肶_j�Z펋k�T+��j*X6*��$�E�2Փ��(?�"�A��Љ|Fe�_�AU��}j���n�~b�`�R�h
�I
�֯�A�l�K�(e���$A�m��K�,L[X��Jj��|���>YOl|�|�os ���ʷ�B�$�m��-`:�U�h��,6W�/�HPU}�ߙ�Lo�ig��w{��6�lR�R������q����]/�}��:x���|��I$7�l�W��ݠ�<Vfd��PU��!e�E�VAD�ߩe)��)}���OG�(_�{��)_V��
a�H$���LY�\{i�m*��;�8���jb�*���K�P!�%_�I�{b�_i��lS����t���Ҕm�I%�?,��c�����{K�m=��c����Sm6Ҕ�����c�wا��m7w��*_$��
�L`�lI$��*�<x{ޞ�q�c�Ov�c_b�{h�l4�k��F6�$�I/Π��m6ǕM�m�^���Ş�m���;���Ҕ�/�R���{ʫ����h�w*��/�=�{c����T���K�XT�h!ZVߕ�;�7�����]6ǻM��=���;��[����Y4S��L�3L!f�A���򵎸�I|�?�̰:����h� D��*/�_/��Pj���1������7��{LY}���i��k|���6�lgOn�=맶<��L8�����������Tذ��v|�	k������E_r����J�$u�b62�YOk�y_�q�[�oR��7���b�m�J�	�/���$m�(u|�V��]�>ĂHk�T�I��V�A��ʠ��A �H}ot�N�qK)O{�{�Ҕ�=�i#�I$�@d�*���Pj���Y���Pj�$,К�*���h��j	/�HK���$�I+T�*_E_�ݟLA#��ë�u�/����K�y�{�{ϙ��)e���᠂�PI)�ˤ\C3 �[d)���^��i�JR��
R����?Zء!U,[[>n���C�LS A���ݪ�I
#`_b��e=�{��/����m���MW�F�ID0A��x�I���2�(A[e�6���}eb��R��nҚ�q��{��N�����/��a��4L`&�H$��}	e3ꐵ�>����TU�W�U��0P8�I|��Y�[]/���~4!R�
��AU�K�y� F�����m����i����D�t�)JYz�A$@$��ï��I%nfY"�T��% ���m��	/�AY]��UPM�$��aZ��}m|n/�A$�_$9�ơBՐ:�U|�@�_��U�~?PE�0�lI�I/ʠ����I�P� ì%Xp�k�P��/�Ay} ����s X����J4�6�(���Ahf61W��P�}�Pn��wGcll����������u��� A���m��%����	/�M��m��qǱ��{�v��2�ǏO�n�t���{�e��N=�n=��/�oz�b�R����LYO{�����q�3�Olx�{o�|__�BJ��� �I"4:��J�2�M�m���%������6[(�?�/��33/Ư��4-vK����;�:x�y�n�)}��pU|�	�-�@��8EN�����ͬ�^��}�,�=���i��D�e��nM��e)S�w�o_q}�K�PL�k���c�_`#̷�W�!��lW�r{�v4�Om6���Y(��m���6�$�*�iW� �[_�Y&�$�E��A���UU�_cc�{i퍴��R�o�����lm�)K)e+Q}�����i��R�YJR�z�ٞ�ow�/����6�����/�{����)B��1�i��cm/ηq����������{������8W�L�lQ_@���C"
/�?5��(�/�1�W�/� �X~X��cO��b��	H�1��ٙh���n�@6��
��_$��d��)�ߥAm}`V�*�,<A%�̐b�ߤ��~6�訛I����Ea��8���i�������m6���}!��H%��r�-�ό���֠Ь>�{c��ާ���{t������ lEK�6����M����;�����/�z;�m�KM}���/�ꂨ*�I|�b�!�)Oi}�yUOOlb��{i�����ҙC$_$��v��F�p�hH!R��q����	�PE`����m2�����w���k��t�c7�m�lm�������l{S�7l!d7E3T�jɩA���$ajc�`�1�{�ޜx���}�{ǃ�B���$4��H%3$�Q�0A�
=}~{�R���������a����T��%��JH�د�s嘳�6.�����m�=æ�{��_M�q�]=����Ll{�P-aU�$��0�eI_���Λi�k���C{�n㧋<�@�j	[^f$��A_ү��cm61�|�ww��4�q��ɽ��?/v6ǷΜ�>z�w�Ŕ�%����--os��Þ1�������6���M�c���OJ�PQ@�R!/���d�I$��������6�)�{���M��;̾Ҕ�=�Ş�c�w�{Ǚ�i�6�lm���b�q�)e�3�\��D��ffL���!B ���|w���;Gb�1}�d���=�p���ا�K)�{�퍴�ATUX+U�*�aV��ka�D�-����:������_}�U������lc:m����tv;��f6;i������|w�lcz��E_*����m�lo`UP�|�T$j�a���+b��5k��0˦
�ʒ������x��m6��6=z{i�i��5|�%m��U�PA�P�� �I/�?TP"�� �_կ���˪KM&�,W&�+�Qi�+'�4�I�I&��$MV�h�GlI$�Z�J��TE&��B��ύ��M�*��R�� v�6) �H��S�������$6�Q$���L��mv��22*����*�aB�]V� �P�5��R�a��I$�KV�CLD�o�Ih���)$�D��m�C!1���[\5Gi�I`� ei4HmMZdr�52H�X���H���I*�Y�5B�l����	��ͲA*D�+4S*���R�a���RI�IHMS-VkRG%v�H0I0��5Yq)e d��K���$�2�B���J���T.[l6I"Aj��>�~��i�%����I�T��mv��I$�I$�I$�K]��$��H�߯̋l?Zd*-���$n��I ��Jd_��-��BV�-� ��h�[~A2��[~����?Ue���?l"�@��m�I��?+l��B0��I)�D��'�m��M��� ��I$�Km�Ih��1fI$���7���XZKB�ZZ���}=�<{̂@'���l?!Y�Y$�I ��㱏xi���=:��o>:R���ON8��ZN��u����JP�)JY�qҔ��
x�������$��$J��$�I$�I(6�UUUUS��M��=��_+�:�K�+�1 �c��8��}^6���7��)�{ʪ�W�Κ`U|�0�?�/�A$1 -��A ���T��_T�H$��|�d�`� �~#0��`�P��� �}Y�ߤ&����E��������������6��g���K<{�{QYnٙ9d�L#MQUMj��T�'v�oʯ��D�
� �T�A���lwt���b��6�����j�I$��-�I$�I$�H�����=�Ӝb���1������,���Pm��_&M�RJ��N_f{����7������8�,��}�{ʯx��������6��m���D0�� �hbAb�b	/�����
-�I$�CB��*'�fG�-/�m��M�6ǽ��lm��;ؔί�A���ݒIEq@�q���i��0o��x���{ۏ�g�=���,���]���m���M��3�lg�S�b�,���d�*@U��*@�~T3g����U}R	��C3�l�$�H/����I(U|�T!�]���b�!�~W��i�6���;�>c:�m��}��������l/{����t�B�%@ A�c�������e��	 *�0q�q|��h[`�Z؂��*���h�
�	�`u��Ul���,_,A��,���U�j�*��;�:oc��R�Ҏ�퍱�R|�"� ���BP���_�_T��b��8��<mwK�m�{��=������o{i�OO{��6�m�@�6�����L��b_,+�� 5|A�P�O�C#�_������ç��<t�4w��S�����O[h��R���H!a,$0f9�5�c|��_cm1�*�w{��=��8�
{�w��M�6Ǻ����O��}j	 ����V��x�&�||P�j��_$�I��AW�;oաm�� �B_T�h%��̒���C��P�}R�$�6�U����I��`A,`���WΠ��$��{��7cm6�N�1B�����EpZ����>�l��*_'�6��0�� ���_Z�
�¢���PT�<S�n��L{�ǳ��=��i퍴_,v6���J{cmi�{�v�lm��t�L}�����`��c�g����)g�6�m=�퍴���m��AWί�A65|�����%�$W�XxF41/�C��$�A[$�k��-��ϥAR���"@�0��ؐH̿Jo@������l�K��S ���@�_$�IG��gʠï�	?�({���<��<qe=����{cl;��1�_{�wy������i��+l�(Jmm�/�PI},�'�_Π�
�`���*���ROm=�w��Llv�)JǼ�=��b�SŔ���{�Uޞ��_�4���QQ	2�0��0���˘��E��@w�W��Z0����'�zc�({.�>��c�?������߯؞�6���4���i�RW�_�o�(8ø���^/���ڣer�Ț��<w���5��㻂);�2��4��r0�4��=��] ���[ףw�����س�Y��l�l�\�\�\ǲ��[m�ý�ڃ�"�3Vu����tTUj��}�9"Omꄗ �0W��}ׅd]:�o�p�Xs�^XEv���e�w�P*�J���t���A�cF��vu���cl�o����M� �fI������aKqt�^��a��.���Xat���'�/����j�ϴH�5T�-�0IC�#U���<���2��c�+ζ����W.��p�.e��K�o`�7Fc�RL����T�`��1M�P�0�F"�r㻝l�+�s{����ܝ!�3s0��"���c>3r5f+�9��9ԝ�7�b�t=ϐٲ="=�̮8��v��6�h��a���&6�����t�:k4%{B�;gZ�V<Cn܋�̽�S��SGT;�	����;��Wcm�iR�����rv�D;��84�7�v���!5,wùtы�d��:U���.-˖)$C\�T�M`׌4��"�sh�˰",�N���4rCp�Y�k�,�@�%4R���/pq�'L��Sa+sS����<r�D9�]+��;�}��Z�A���vܝ�pǤ��YɅŹ��a���<�/����\6�������H�M�}Y���Y�w8���&)i�ov^{њw{~���f=!s4�E�)p7m�~��GHn�=��Y��uTq97e����vevq6>ަ�Ur��&��mj���dyb3.�ܡ�����v0�����wf�����%��WLم�b�G1]�{��vE_�>���>�v�飘ٺ�o�.)�w+a���0,�%��(oY�}a!Á)���x�ݭf�"�~�{.gr�1�p��c*���i+t�e�4��;�;���Q֥`��s7_f��7%Vl�;���ǿA�wf����X�d��5�էq��G���
+x��׻�wF�sg����k��M��m0Y5׮Isu�A���J��n�׋�-fnfM��I�y���%	��5��Y7%�*=��ũoOj�|��z�j]�k���p�ʘ��]�q���J��r��8k�R۲q�i���>��>Y>]d��=l�-R���
���KϷ�l?{��)�G�^�	(�zQ��$�s�n����h�f`���b�`薀zI�s�{�}����n�#�q�n*K;����Gv���-�!tN��_NW�-iD������5�=XZu��n��m��8�+{��4l�h&E�"l�H�`�09�.�NB��RѼk�R6齑���C�6�w�7�v�.+w�9.:�P�,9�3���֍��0��Z�f����1��n�LLI�9;��	�;�woh��s�弒�[�D��\�c� ��F�-��,7ⶽɻgr�1^�fkkYf���.�֊Uɣ&���J� �����uh<U;��<f�][:dw�:n�d�\ow�\���7�EkwV��K��0�Z�x����#����'3נBǺ#}4o|V�Nv��qs��應#7%� ϻ׎���FNz_�嵼K&js��32��y�v̖�����)�������=�d��2��{�\tΎ�����}n�V�L�8[��M�^M�;���z�'i��|6%D���鐪�zU:��y`h�2�[s�h��������M�8�~�K�7���X-[ ��U{6#H��tmh�R;$3�� �*x���%΃h����
�ŗ�'3��P��N�6߳w]�wڧNww7fnH����G^R����|����7��m����\�
Zk�=๰�-��!�����SZp�&,m��2$�Ah������f�du}�nظ��[G`"=����m��]��bS.fr˷&��'&�"�W�wv��\��31q���.�1	������V�1�Κ��"��9��̧˜�A�}�0�F���@噭f(�Q����ղ�j�͂�//j֫ed�j��]�\�	�.��=fŀ���*���q�}����r�x�#`�%c}��|�^i\�nc��Q���Q`�f��^Q�BZ�i���P3�wJ{^)���M������ݻ7y���[��F68�[�鈞=ֱjV�j�^^3��7W6���*��ff,�1ymV�neY.�GG���D�؈��h��qM��fw�ʹwr�f�Ѥ�r���K&�r���f�J1tw=\w���Z�%���a��QY�5��L��H0C�0��qݲa�[Ĳ^sA��s�S��l�2r��G`�s����J`��Tw�e�
�_��b�J�W#�'ps:��c�l������\��1m������::���-��GfE�]s�r�C����K�(��7�K�M��IF���b��6m��Ƶn$6NZ�=����6���`G�F:W�,�M�ؔpBC!��΃��+!��9�Fe�(���$��k�k�]e|���{%Ӈ�Q\$��q�]�t[	��t=�.���7�<��M]H8�c�@�3�ί^t=�M�q�3FMy�	�ϖ��ՊH�4�)�{ v�{-@�ǎ�(��C�t�[8���wټ���"ᮾ�y��{�1K��\��+mKrML�U[Z�+w8[�ܥ�E��^�d��\
���n�)?=��/p����f�|�n5���Ӧ�j.K�ek�0�h��UV��K����_��b]7�iuK�M_��$�z��ۜǹu�z}��C����$�t�X��=���50-�r�J,�>:��SeC�����x7��o-��������L�7'�N�yp
����Q]u��"2+�a�F��s���Ů�Z��F�	⬒cQBӒ8dP)f#"16�Q�dR)$m�RH�F��h�b�Z"�m��Ҽ�vʼ��*��^���m��A^mtW���*������l������]U�j&(�ElH�h��2�BId�I��H��l�I#m�a��#��HKU]kֽ��kNu��6"#�!r1FDI2C$jI2!$�I"���^UUQUUm\��$��Ԉ�R�"X�C"��I$��ڂ6��lUUV��U�⍮����jZ�uuDWl��{��m������gQmUZ�#m�mkz�m�Pj��ʨ���W��[U5�.��b-]��Vm�QvȪ�����j��l���kZ�h�-^ٓ� D(�0�&F�0BD,6#i($�a�$��ȡiF�H�#.F�׭��1��UTm`H�FB�.�qC"J	$��r�?72"d���R|dr(H�FbrHےI$D��D��$�L��KiJB%BJPI�#�$$&	$�G�$��܅��2E	-����m��������kj��28L�����%1��/�$H��Dd�Bd&	$�(�QB�e�	��$�I$�AO�Q�nS�n�TZ�m����G+h.L"Z9$�FۑH��9$r#������m������4E��sֶ׹U��W�5ms`�	�F�rH$0��$�	�$��HI����I$�	��RI$�)�����[ͯ��S�k���P����a2Hd�H�1�
$���FY$������$�b&C"�@��kmmsW6����5�-���5UU[DiW\����UU��F��[V���-��[l�{[k�7^3��UF��k[\�E��[U�UͶ�7W�z��*����m���)D�I$��Hܒ72��	#�I",'�E$��M��J�ƙqFL��	24LfHɄC	$����(ڒI$�H�$�$I$����	$p�#$���$n|�L������V�m�m�*����!1!	dȚfd���	$�ai�!iL�H!$�$p�F&�18�P�"�Eq�$�I? ��L2G��%�$�IP	�H�km�ge���mU����ۣf4$P�q��%"*J�D$���-�ʪ�5WF�g�mE�/aU���sv���km�щ��&C	RH܇�0��D���d��0��#hG!$��I$�I$�6���	3��d��a���q5�UUy�����6���m��Q��*��˛im@�$�p�I$�P����nI$�I#�(dD��C&)��$�dd�ܑ�Id�#q($��$$�ڈ��$�#rH�I�$���\*�j���m��m�D�$�I$�#�L�$�1)�U{u���]׻�UUUUVI!2I$�I$�"$�قH�&C���2��C"p�I�I$��	"��e0�̑%>�CABI�m�����UZ�����m	F$���"�9	��Y�,�Id��$�L�	$F)	�	��ko^��u�6��m���zѵU[U˘�������o]�6�a��ں��*���m��˗5�k�����D�$rE"*#	�I$�H��I$sv�u�j���۝UX����>�Zr2R(H܈�	2G��nI$��$p�I"I$&�1�HL���F��(I$�Q���A��lF9�7	�	!��$2Q捫�{���r�U�)k���]b�ڶ��xm��][u��u�F�ֵ�m��\�=UmF�v�\��W��ƒ�F��9$�FےI$�H�"���pȡ�R(�1���kF�U]��j�m���6����{d��*�m��α�s[mkk�EUUvm\�ъ�*����k\�m�"L�6�2FH�A$�C$bERG�e��$��A$p�Q�$�H��݁�vW�y�m簙3m�m�k��j�UU{�h�jf�ͪ�����z��In	 �T2 !�I�	V�m�Zۨ�+���k]\֊q&I2G��I"e� �	��	%��D�$�A	��a$�	���EUj�r���oZ�6a1H���d��"(�$��a*HԊ��>�FK��$�.G�˕Uy�j�E�m�d⊨�sZ���k]x�k��Z����Yo-����^��溋M^�j#��#���j�5��3�y�Wv�dW5�V�s�mUQU�G$P�#n2C%�d�Ha��	-W�W������r��b5�S�r�]kW.\6�xu��Fض��������u��ym�QUUm`���^6�m��km��m�݇��Z���W����2Ͷ�m��m��m���m��m��N�-�cV�EUV�Z��ͼ�ޢw=m8���[M�m��Z���P�䄥!��"Bdp�d2GEy�k��u��-�
���h��UU]��*���ڂHɍ��rA$�I$���^�U]��km��m���m��" ���uU@W.u���m���W���"�6�IH�C$rI �InI$����df	��RI$�IR(ڟJ�m�UU�ov�"ڶ��2k�a&I���H�R)$�I%��׻-����nUUEUrK$��I!"b��j��Q.##�I$�H$�Y%I$�2Z�6䑶䌶���&H�D�a�II$����S]&	"*"I&����C"m�LP��I	��b2V�z���C�U��m�mv�Y$�(Ʉ������lH�$��j#�UUA�ժ�HOů��I�!"��RH�jAaRE"��I$��%��6ᄣ#�%(�H��([rI$E����]]c\�UV��ͽAE�UyA���u�ѵUE�[���kUUUu��u���.)�I_BL&䑲[Lq� �dR!
q�Rf$R!1#m$�I
$�#��H�%a�<������������ꘫ�ەm��]V�V6�$�Y%	FI$�O���$�B�D�I1#���&�2G$p�Mj�گ+�<�5W��m��x�H��h�6��*�mv�	2DY��$2I$�Ha29$��$��m�$ndQ�K0ȡ�DQ�	$�\��EFЂ#�H�&,�Wn��v�5^W����mm�b�um�W��^:ӎd�Ce ܒ&I�C�

9$�I$�H�iȔ&H�RG�h����my�UW5�1m���+֭�������eUUUUm��n^�\ֈm�UUUU�.��yrڍW�T�u�ET\�{�ͨrFۆ"H��1$nH�1dssd�9��cٌ)�Ѷ3��:X����d�Hlrٳv̩-�� D
�o���z�	��D0�����ѯ[l��@k2�OB���
~��ğ�**�0��*k��n������������������n��n�n����V�f�6����n�<�������l�2�Jޭ��f����������������W����t5a�Dn+�\^쬫��G��yzL٣W�<�C�D���O`U�~���Vd����r��r�k:��]M4��뼭����56L��Z��՚�qm{q�ֵ�E)Ux�S���\�~���V��ҭ�<�<ec�j�df��K]��g�w��շYu������-�25YwpZ�Tr.ܷ�&��Z!���V���[�|M=evy�<�t�9�z����WL��Gٛb�þd��n�=�s�\��,�����N$`�T��u$l���5q�k�U�h��3�N.�׺��a����7�6vf]([T{���FG�"A�=U�Мf��/K���r�<!��;��{����X��1�c�K�nv��诒��z�O.E.��:��d�w���N�������Nϵ�����͗��S��wU9��f�Wa���3w;1篖�fU�{��wǦ��o��tiy<��z4��<�]�������C������f��Y�����x��٬��u�-��ln8�V˅�3ޗ�4�OfJ�:F	S�4;f����nl�1N��S����I�nvygW�4x.�Y�Y����ن�m���]�My���d��\�\<�c�c{��/\��\�yl��*�*��m�ՙj�f쒞%��x���L�CK�����=�ao>R�:���n�ϓ��ʭF��^�T4�R[h�C����9�Xc����F<t?3�w3UZ����p�.�ر�H�1��3�a;�w���e��;iP�n�L���*���y��9s9t��>9-+�="沪ʴ��#J���q�S�9�J{�����k�k�CR�ƭ=\lNN.�LS�F[�B��,���ʭ���f%��<�3�N.k���Z�u�14ʱ����W�u�;�V�Q�����ճc�@ՙ���C[Ce��Mv�f����Ooo�bb����2f�ų��{R�y�]�m�Ե���w���]�!��j�n�Yt���^��fk�l�g�؜Ŷ̅1��Y�e��ve�3b�Wd�ڍ�ʍ���g*�/n.����}��r2"�֔���-��1'�ǈ{سs�A<ٲ�fZ.^�V�ؘ�v��.u��ftSu�.E����1����h]�����^�s����p�]E���{Z��z�3s+Y,����&=�Z^95�/��5�m�/����O������׃˹�^�<��UֻN�-���;��+2ff��B��L����NMFNe6�ՓyH�y*f����+�9���m����t��R�	����-L�de��K���Ay:��mA��^�]�9����.c���8���;�ި�c���^ܺ̽�Vb�ĻeT5���M35O����eM�ͽZ���m�/g�#4����>�v�>�sx^=r��nk�9#�fV>�ʹ�^E4����ʬ���œU�Z?q^,�XU\�f�x
}8��7��SQ�ٕ�Y�+�[����v�mu�nTY�:MN�,:�:��9��+,��}�cy��s��ӷ���g�G����Je���t�x��i]��������'t�h ���*�y>)K�qx��v�t�`�1`�U�j��s]ۊ]X�.[Y��z��b�'�g�+��j��L�$|)�3V`��4{<�"�\�Q�y��Onn�v.f�ݎw�4f��9N���KX�\��u��������O��$�ΕsRC1�*����6L�xm��th�xy�k93Z��[&mCR�J4Q6=��[����yf>h�x���df�oz|i�=ё�\"z��/:�|�T���-�
K��0��b�ɽ�
φV���I�j��Yٲ�U���,�٫k��R��t�2{�P�]_�q
|�QKEֺ��MME�-S�fd*����M�иr�Eu��dS�2��i=���w�yG�MMW��տr�%ȡ
%m�j�d�q9�]o��1f��j)�n�FV�-B����95u|�l
�zͯ+q7�{���底��:�ra�r��N>�3d�K�V;��"��&��^RR���vZ�{���`�y3r�Y��"oY�ֲu���Yn1٢�wa�j��'b���6��seiI��|I������]��j̚�g��d�5�;�z:��c�4��Lֹ�y;w{���՘��k��nF5��u���IQ8˘���#3Σٗ��ʪ�J�5�km�6U2��\�I;�>��V��9��^�[μ���6N��^`�뾝��õ.}}��!�G�L\���t�����W�ޘ��0o�/{������h֛��zZ�˭+#E\k�ʭu-����w*��7ȥ%��b)Jg��Ǹ�Q;����1�OC�:a��&Ė6t�X+g-wV#v�Y�.&�j^5f7U�i�ڪ�z�i�Ŧu�qi�X�˸]�z�Ǘ��\�3R�6rU�V&�6�	��T��xu��-�U�lY�jՒv����vŝ����,��5m�^*^Zɸ��Y�-2�M���y}���n���sHS2u�t�z��x�J���t�')�\��YVT����e�G&bg���o���_H.��M����U|�3-�w�]k�Z���i�qVq�۵�*�b(\����k2]�r��'5�����w���E�5�����OR�q⽋=:�&���@��NzG�D����n(7���!3�1���_n:�5֨�\m�'i������$��m�0�ͧ��֍�66��Z7gI}����m��2c.7`gچwi|U��[}.�w"�zاRp{sm�W1��2�/.�
f�#\f�ݢ��]pmk�2b�iu��WWlۙm�|���Y���C!�<8z{��n/4}2T�F�]��L�ek�5\�=�ܺ�ދ��wy�^�S�����nR���\��[��eFK^�l���i���:����Fd�kEB����wOk���Db��ٹO�6.mR�c,�-��5���U��cnٙ���>��e�(�3Ks�Sd�h��7y�4Un��m���[�=ln�i*�5y������V��n�|���;�0��N0��VK�<���'ċ�PEF�r�Y9Nt�NO���8�	F����-��p��9�͢�1eˠ���}3,�6	B@-�dg5r5�lVu�x�����/ܧ��Z��A@��
S���?�C����P�e�Ot����Ŗ��Е-l��)lY)Q��[�`罔>mCM	~�y����//�>;��쫬^/Ls���z���]�b�Vr�[o]^sI�.�5f��xrjBHiS-gG�T#��d��y]�쏨��s�]E$ɬL�!"Վ5����������õ�	8�.YV���^㞇|���{>J��d��fT���5+�8�O�w��[�5��"��L�o����;�����q�պ�"���ʲ2�R�7e^"��!oeV�3g"��z)i_j�e�ʥ�܌������݌33cK��e��ٶ}�,�OI��}k���Jk��8��˷���	�v^�j�eUVi��r]n-۸�aAF�;�T�}<��f�q8"x�ޞw;���9�6T�2μ�F��Z�`S)�=0�˷7���,0c��T0�̒��>�e�m�u����~E����J�Ȥ����������h��`Ȧ�֦N���hT���2��Gvqs՞,r��I�	�Z���҃m�=z;}�%٠�7횇��=������;2A,ˮ۬U2̢�@�)u��{�������ᘸ�ُ�-��P�yL[DDm6ᯒ�
��QTk��l�o�R�q�����1��=t����ػ����3��zEd�+NT��R�n��f�dd~C`�X"�wǦKܔe;�c�]^��#��/)7�.�PZ��X�H3�7���&� ��<C��7ސ�i�@[2�PSť:E�cv̙�bn.�Z�1�^�Ƹ|[g"�Z�w3f�.~�߄Q�p�9H*�f)�qG���#����vm�.���e�ҮݕfԛdkNd6L�O�3�(ڻ�1;;�ón���W�:�P]�]QB����UK����o-�����{WW�����n������;T]J�1��9V��H� �nn� B%����8��]�|}��� �R"�O�}�6��u�>5neiw7�>����橴[]D��樸�g�m�#��]$Vu�E�g%7qA.ꝙ�L�b7"Y4i���֕�\y;�v���q4z��:ս�1z�ъ�~�PR��v'�`~�h➉��c�K>=���}{wN&���(�a��#Y�6��!Zw�r�pȗj�}w&&��r���fw"�u���{xz�i��.ڝ�0ղ3���)-]b��l�D�#�$�~���}F��¡��Fw�מ�b��},�n��-��/2�ٯb-V��e�s��^��X��e�{��W34�X��V���gb��p���q~���O�{	㏟��A���Ǜ-�<7��8�K�l��A�p<ZG��Њ#�k�2ۦN��{�e�k)V�e�.�Ի�D�;T���U`�r��:�cc��^pͯ�fzeL)u���u������R��-Z���o���Ш������}Y���{�����-��V.>W���o܃����L������y�A.
Onp���^���e��^v���ǖ��bBV�6�<���*3����u��n��S�W�Reˏ
N:��heb�\��M3<nvr[WȖHI�aI����{]P���b�H����ȳ��k��w�5O�s��3�H:|�wg��V�瑌ɛ�[H�s�0�d�p��T7�x��u��&����b�~��w�i�#��W⋽֏a�ɼjx������M��}ek��U�4�W�bV�9�X�Q\c]�b�������Jm.��P�yt���;Wy8f���ۥL��V�d엱�;�
�2��vd{ڊ�^n�X�l�n/nl����֟W���\��$�x�Y"����eb9�!�qc�^9�o�/�A�k1:ڱ{t\�L�9��ň���:L�u.9y'����hy�R��1>�t���NW��V���ds͒P��d��%{[�G;F��*��S×OU��Mr�_ov�Э	V�:`ә���Y�t·@n�|��ҔW�Ob��{۝I��3�D��wl���<&nwl��||a�Y�7�YK��V}�)׳�}2�s2���t�^�N��Fm��Wl�zL�����[�X0�����3�_��ۧ0Me����0r�V��'{7��3����v����y�ot�n�uNP�x�ת'0'Yt��ո&�GQ�i�񰍸Ձ�j1�d�-��q���f*��a|D9��e�����KB��(r*�v���y�]�e����P�kf�#Mv\K4�Γa9���k��4�Q*�+�O���0բ:�8��]�n�k����:'�c˹4���b�f���ͫ'e�d'_f��n�7b�w�b�g3����ڐ�0u�#��=,�����;���ΡU�����*{��Z� #*w��Z���������\V�6cS�r��*���Y�Y���m�����f���BB+�
�p����6��fwwU�������an8`hztۊ�Vn���v�D�8�s̮kښ���X'�vC�,]:wO��<{�,k����1��1˄ �3a�v��m�(�	%f��uz���m+��v-�.fz�\&Ӽ�s��F�1m��b�x>�=f���B��X�
���M�\��;^=���U��\;��
Ķd}���I�e�Js�սV�*�^>��OL�<g6`Ε4xK�س�e��~�%,�5�-��yM�{�n��Kw��
�,ۊ$'��n�C.�����VG	��K���e.b\�r���3[8J��w�z���:��v�qŵ��W�,Ä�s�p��Qjϑ8Y5Wc�C.��E��*��]�a�pix5_�y�J�������,2����c]2���>k��K����f�ķ/�E�Ř��-N٬��cW�<��#�𙴼��hb���RV^�����kے�o.��n�g},�l}`�l��l֒N9�9 z��x�W$�K{�wk�>"�w6�M�'��6M��u��E"t�2&V��\U�fen��n�������m�6�&Y&�U'[�{w�2�W��B/M-n�T$6�{u��)��9�DPHh�<^: ��ky�U���ETz�ѱ{6�qR��6F�p�/n� 6j�ge��6ҭ���-Tok`�n6�B�� ܎O� ��-��F�a���l���dA��D��"6�G5W�j���e����E�aۗ����ȵ��Z�׫4UPA��!F�Jl�wd�Xu���]Ʈ-��da��4�(� �x��S�O�βOiX��Z#�'wr�4WJ#\�p�����k#+�z\�Z�wKܔ��l-�lķ�UH�QьiX݄�WrsɅ<�<��N�������Ŵ[X)���Q��-�gB��N4�v�T�1ͨ��3���h�ʶ�9���{��*4n�G��ãk�f���5���^�l�u�j#�^Vce9�Q8eAUH�UPbAUb-���α�Ula�!H�g�"JCJ6܉#�"�6+�8hD�f��F��y�[6.�4uR ��y��4��*�kFі���tf8sA��<�X-�dU�װ�y*w?v0��D������o5�w#$:�@Ӎ� r(�f!$�ת�X"MD�X[j��"���]u�k�r���+"�^b"b'#9UMD^�ݖ�ɝJ�U��ʼ�G9sZ��s�"`b0��9/e^j)]Xփ`�F��{\]�m���3X��`��a2��Fʋ\�5�`���a��:4��3[h����"�W�Z�"�5���uܶ�du��Tr�9���Tș�z�7���5u�L1�7���Ө6T-���m�*��&N��K���E����,�i[U\��/5��*����MQ��V�����ΰ��Z�9�*�n�9+j�]VѶ:�N�A�h�;���m��{T�XTc�{��^�C�\��:�f*-�Mm�s���l������r�"f�{e��ײ4Ơѡ�꫖�^%8�Te���^�ݐ��mE	]V�vȥ�Wf����ʧp5{NkJ�uN��͍��um#l\c�C��"-�;d�\�ؼ�xLӆ���.�lDݓ.i�ƹyp��Ey�]���Ȏy�u�ys�PG��ǫr0�@�p�"�����m�i�l�"ڏ�~ߟ��pF���,��On����>��*׳��^kZ국��nz��]��ｳ7��+4�n��r�T{̗��s��cgu�'eU�V����.��/m^�;d��;���>²_{ب�5�_�A��*�M{FyԎ�0�������jyH�u`�/�z�;�/��Y���r˞U�y"�Q�f��tY�wl&1�f�����i�H�k�cw�v�����O\��Wu�}�q�0r�;޵,B�o^�=f*�;i[n>�*�+4γ<ccĕyNI�QimL�v�v~��L�ċR-��op8���Y���a�[�{0k���7XUݶ������|��4�嵬�fb-w�:��q-����MG�&�R�J�*��목-zNRP��oͽ.�ݍiv���l`�غjiii�5�z�q��hn�ITQ���뫁*��.�)���������1�<0�k�DS�"""�11�ƕcD�[z�<��������㦝X//43�Q� �EQGl	����T:m��n;��p6��Oy��ڋ ��"!�Ra1�t�5Xp�r�{v��=Z�r�X�'(�y3���N��b��G9�Ç/qL=y�R�-s�Z�����"�c[��Ny9�ңvy�����UV&�<�)�Y�^qsm�)Yr�O���D��ֳ�}�R�8�dl�]�*�H�r�8�~zk�{v���/nװa�ױ��Pp���(��I�o�b�g�C�L��K�DrȐKAv]���c:���D��B�h�����a��s��[�ב���z�PW/X@cz�$��v~�"�������L,a�qHF��Fna�����@�je[y�u�~D}��t/�]�@���$��G�l�2j�m̢g���R
<�̉�����JKK�ҁ(lUOۨ��\��!D�b#b������ֽ{yL��%�lDաu�"GStH��4�߇���|L:92�K�9ɪa!������ U
(�_E�(�]1Ч�����a����d�OX�x�*��*{D����j훖��3H6*y熂x�D�Upq�Lq)	���Ei��U�35���3L��2^&[V-�\|�wۺ)�W���Z�-_b�e_^�cw([�ͻx'v�fc4�{�lȅ�|����ZX�X@��j�ǭ�gΚ��50p�~!B�E1Bҥ��"�v�Q)�c{-�����W�L��%B�S="��m���頇/W+���1�r���5�1FP2��|�jڡ�U�5i��0)ԂH	�筳���{6#�u�*����dNt����;�sI�Ӈ��X�32gG8s5c�m�����9�s��hN!�3���)VȁЂ�tL��h8��`�q�dZ�jV����ʰ%qi�8¥$I$�P���VBq^��z"�.:���p|Z����*�qn��.�8$twGB��Bc^'A���`��{�Z�^�j\��I�Uv�r��svɑ�_6ئ���cc-��v��L�ʼ��םgqv�I��}61����9�g�A�q��̊�K�q�$r1e
���s����CW��1��:D'L���{1�Wi:�0��I$�A�C�����nTNJݚ�T7_�l�"�)���͕Gg�^%�-rg93�/S�1
w��>�>|�΃�������w8 ��`�笷I,��2$Y	Hb-P�눘Dg�'�,9a��1Z��$&���hp%�(,ҝ�E�F%��4Ş���v귰�C�ܶ"z)Q��#%����ʙ���񥐻T�� a�uXi�Q~��L�Z�b�k�kq;P0Wt� w��!r �n{��b3�rs�L�j���Vz9G��2'uU��傞u�miY��l�ʫb���^iچm�j�-�Ƨg����v�}��X��h}Ȭg.���X\[�y��r�ȠZʌ4΄��$�:��ib���Wmw2��î���1������8nXhhhh�uh��E�	��	�.���Fi�TP(��9ɝ��ሞ����Ï�1b:@�gB�B��9[�򅠔��B�3��ưm5�IL�A�.::a!�!�um�D��7l�Cii��:��o"���֡�3�
���μn�Jp	G�9(�#�ۈ�ш�o/m}wj��n�>[�H��B! baP��$B	���Q1�5��t�\�s�� 3:s��4�S�ػ,U�i��0�Ar�x���(C�[�KrMf�h�d;�"�FL����m�������ٜ궱&�'Fj%PZ�TA�ƻ�m�MZ��3��35����9\�\��U���\�ʪ"��l��j���=�}�?����RW�������ͅ�M�t��5�Ժ�K*��D�ix��0�ұ�VTL �\��j�:����qU�p<��p��yU^j"�WA���z����N����s�;��<�i%(�]���&:���c^��K�2k"/=8�q*6���
��6������)޶\u��®V^_o�z�ڦ�����;�
���'�W;��MR����&����4s��s�d�A����5����D
���$?���'͋�ۻl�r��E��K��d����4h1"%��@D*�����VH��)5L�:���(Q��E��,�BF�Z�;��{��� �#����B%��`�A��$)T
&J�����.�fG.�˂��)�w��hr1H�-�FW/=\_;*6C��%\����b!����RԶoV���0�{�i	�$ A'Bu�!�OH*�ˉ}/�{�x0T-:��������M�2���:|�$Z�9�a�	2���27�ߟ�_��O}��tL��^�3�
(�0X!�
�޹�w>�Xē�Nf��.�V/0_W� �R�i��s;��R&A�93x-�oLgT���q� H��)�7dV�H���z�]����^m�鷪�̍���]�5�X�m{�Z�hli��4x���zy���� ��t��a�[rwBv��@���B��X�L���\}&E{�U�g:��9,�BIĂFc�޺TNP�P��K���ǥ�Ci�W��P��'e���0Ⓡ!HDx���u�ڗ�z��cyQ# �}��{�#�&k��|j�שԡ�A�&I­@'�ֹۢ��j�x@k�v����.��J|>�9�^��s�5M�"Y���qG��s��8ta�&ƜS�1?_χ��1���ސ'H�6v�.�aj��z�w�cj$6	S����F@d�V5Ñx^Z�e������Au��G��#�JB�wdnլ;�&�ח��,�HH&E@�2��U����D,"�kNb�F��|t z�o*����}��5��j�VQ��S�\n.elM2��ۭ˙�o{q���֮����6��P�f�V�$DD����D$"C@��͢�t��UGI=Y�6�)PՈ
���o[��6���pAie9d<���aJ�"8�/o�r����=}�>�����x#8����}�9��s�k �2:�1?{��������ߦ�����s�L�:"C���M
RBA ȑ�܆���CGa�t�r:��=�=|��-�@ܲ'n�&���rI$$����;y�d\	́Y�%c���5s�;� �&�c��$���ʙ��G\Z����)HX�9�"A�����Rq�Q���ql�=����T�V<@��C���f::@IK�R�f�,!�B=W�P�È��ZF�K��ve�,<[�6I�+��N�3�l\ݭ�dl5����L��m5�Vfn%ix��,��5A�α�ﶪ��[��D� ۑ0XL����JI �'0�\���tZ���D:�s�O2���s�����r��\��i�B���d�p��u-5`�F^���'���&�g��s��8��#WkjF�[ �!!����]Pa��v�ڧ������`@b�\��9$��q�D������:f�ّoy�32�/ �1a�����*���d�|D��%%�t0�R�uDe��b\L���d[�h����ŜM"P���Iʾ��f(G) �`���A�'^'U��c���)$G�P���Ph�A�q�����i
�L�A��B! �drM{@�j��[;��#T2vʹG�|�}��|�ݧQ���F�R�)lb1DaD2t-h�6:ĂH�s����9�ñ��7<��׽����޺z�Q��txh�Ȉ�
�dUD[^*G���\��9z ��&#�D��ߖQ���'���[E��SX2em+��c��6b���b	 FF��ĩQ0��ɓ&�QH҆#����IV@u�]U/=�h*��Nfs��*�2I#��p�(�7!�Hѝ4�k��h�瑼�[h�ӕE�`r�9�Ƃn�ᐶtއ̫�Ƨm"m^���&�i�v��;�C��|>a��TQD���(��_D4c��s���0Ξ�09Mu���{����丹��9,#)]؞ɎA@���hr �i�Aתi�gj�gU%���M����Vd�Q�`w�������"A�^�4M�d`�vܝ���)T�$I ttr ��T)�P3u�o4��0~�܈�Z�DhsvP�\\Zb�t*
�F�1�7'���fu���leD��R��ȗ�����D6ۻ4��F8r	���Då`C��q�zN;��?q-
��H/���OQ�]��HrgX�3�:� ��W�<m�P��(��B�(��(�S6q�"=x����}��1�E `�\���\ȱT�켧A �i��s/V*�q�K~�d�D}BHH!QA�c&���mZ��5���{uj�����2�ۍ!)�Cu����[.vn���f�-�S0�uVѱ���ͮ^fk���0�+ˌ�*Jv�	q��Ze�]γV�" �;���CB�W(F��
��8�1}GM-ud�N��V��� Lc* �	e�" ��\�b-L���$"K_L�#_e����֓˵��n���N�����D!@�(��(���SKv�����W.���t�Q\�%�#�%��WQ��B��A���� &�_���?�|�s�����L�1�ቖ�&��A�HHDQ*BW��z����`���"v��y�u��D��Ӊ�t���,Ӂ������u��S�z7&�����۶B$�:�zf罛�ʝ�ǉ$�
pq- ��
Z��y��@���@�	�ә�w~t�-<���=
��,�d���l�ľ��"�}�'P�0�l/s�;�q�}�N��B���Y_��l��i8<�=�32ky�d���PӘ7^7M׹5��щ����=®l��K^�dOf9se���K_Z�)%25���&E[슬�;<N���ɥ���Y����<� Vl鴙���)�3ͻw�!^�H�x�ܼ�ڍ���g%G���zwz�]ʵ��w[�������1暆��Zr��=���U�f̖�	%[��,3MN2��n���~��QWS�_:��������~��mW}��{ٖ���]��F�[{��5�.^bȦ�4iyښz���]\�q�1�s)��\�'x�d>VS�TM>��&*��6���i�o'nubՅ{��\w2"V�-�����Y�!�c�]P��5_pξ���Lu;:���y���WEMH�{,D��y��R�qm��-T,�J5��RW���
qov�Z^�c��A=8����w�l������D��,^ui�4������]FQMwR�W�C,���l��ۇ��{!1s���Istlݽ�eZª��tص���Dk^[�M�>�j��l��\3�C�E�+�3���6�K��i����s�=�n����pm\�+���N��ҭ�����q���|�<G���9+���]�,wۮ��BБ�]W��{��YB���UG��UJQ���$�V�T�IVZJ�R�m�nYdE�#t���`�����#&;nYw�m�ǫ�Z�"Z�Kl���A�6��[�2 �|Ҷ
 �����I��n�
ޯ�C�~�BA	4
����#*O�㶷�����%j-C�
MB��ӛ�A�Y%�O5���|����&�n��m��}	T�x�:�����~VB���~j��L��KS��ip�����L��sϾ]BA~�A�TUDQ�%�+��]/h|B�~Z�&g�QgN�.L�1:��g2a�0���������8s����4���!
"�'���ah�9o�t����O�"�y��rr�����*���U�A�����{ڕ�j����׈>��lHeA������Q$���q`bGP��GTq	 ������T<K	\�ȄKr�����6�9g�X����B��Y׆��mh����JY�H����.&��r'�"s�׺�Г3�[TF����o2' ��ݩn��I��$�ȟKX8�����QC��$�8�!@J!��k�s��qW��
������#	Qk�BT�A��*�� n���"}>������I�
�����n���1�Y.CV�l�[�n��K����z�YY�R�Y�����w����-��=��r"� �zy���\�<n�<`ɭȒ���E����9�.8S�
��̽��g_$�Q�NL�v�Ԧ�����&i�bk�>����޲�G9��Phd�#��8�Y��@�0:&t�9�pL����0SǛ���-��M5�R��aK>�r{����6����D%DuXd4E�}y[��۽f(�����52/��j#X�wsH%lpɓ&rCq6��Z���C;��[=��$�o[G�"I{
�PO�Obf��AC��kt>��B}�O�^�%��TAC[�88�$&�L`48�n>��
�!�K�lGW1�QZY���쾘�H^_(��*��&`�}H�%Ï�=�<����	����*����pQ=Pbg�^�RW,{>����n��+�"�����,!��ei3�1��kL�V����.��ˀ2E�2c�1����m"��_A1�;�*��1O{���܃����D�""� |M˗�OK��')r{"Wԡ�/���Ǥ�{r�i*�v4`ã$����RR���1k5YJ6f�{j��D:ǬΉ��������ZT��D�T9� ��TF�f&ڱ��1�w<����'*G�ѓӯ��;�W�|����ał��^�6�m��i��fb�һ�A��'�1��A"4���rgc8Jk�j4���r�A�s�G9��'�NUU�'=0�ElI�F��9��y�7<��rq�婗�M1���&��:4[×��sUܧG$`E>@��M�$B��1�w;=�/v"�Yn�WU�f����M}����Q4�~�Ѣa�s�fL�c8J2lZ�i�0�s��Ó��	$�Xj�ۤK%)0� �T$3�j#����]Vb�o�\����I�,���y�$�Ug^��⭡� �������}Խ���g\ c�����x�a�+?_�!#k1����_;	k����	d�����K&bW+@HA1�׭Y�f�c�6�ZL���R�	��R�a��W�]�f�����`���D�, �־Q^]����N�Nz`HAi@�(�X�W ��7pYu�cO$�HH8(P���d��5z;�>�V��dO�n�L�[��ǾW+�1p�_$�I.���w'��[L�h'�eT(�Tȃ��0rF��P$)�P8�tG�A��Iƀ`T������W{��9�4Arz�:��J�Ĺ�i ��k�A��|���ɘi�L��L��h�a`�	�;��s���A3���4��ڈ0+���烧����L	�J���:D>���.��שZ���䨸w�!�>��ɿw����W���@d�$���1pK^<�2�O�$��(p���z��8R�<��jq1�]z�U�ƪ-}=�J�m[�������AY����ٻ�P��C�^&l�mK�;�FL.;�]ij��دy󃷪�����ꥭj�3�п�^&%I�E7pL�@hOVB�{�����[�v�@c�4�@���^Q!@��M��ה2;]���Rn�,(Cܽv��MQE��QcZ�B�fVB��NN;��
�dC+�`���X,��:��LG�=�<�*o�!虖]��C�Z�~q_�'�������g���8/lڷ*�pK0t�v[��a�e>>dB������k�����Gf�es2�����X���;�RA�j.e�P%EN@5�*�-C���V�s��[�ɝQ�^�?�'7�>g9�&��s��6t�f1�鱈@�F�X�QC��ss�5҉ެA��h��E+UP���'��W��=�+��x	XC�p�/Y -�P�L���BݳO'xq�L`����;��MLAl`���ɮ��\�I�Vh��{3�;z����=R\C�K=��側�b�q�Mv��y~�W�M��aɇ��u"�n��)Ϫ�{�?b�zWiMÕ��e���]H��z'e�Y�^�r`hZ�Yg�ۼ��1i�a�S3rfq�+-wV��vc7�z\6vk1nʬ��J�_NV�����&"�!�b\�[Ƶ�
��!��Jq�!$��)e@���׵���9�} �&���5�GLE3����zq6�51��C��E�i��y��T{̃*��j�'�H2I�RI5О�NS�	Z^�0J�*��s��%c�s��q"n��Pr�"��-�zb��3h}7�L���؆$��@���?����8s��(�/�@H��矎B��`"a3��9�M��g8x�Q��7(0��J(B�U@�Tcr�4���De����`6AmB�v!h��Dz��z}�}�Խ�'4���=Jg�� ��˲�&@H�(B���J�HR;ձQλG_P�I���R��I�
�nĬz�e{�@b@��O.�Y�%�U"�;8th(�f��4�	�Q��{t�Z��k��ow����/����{���VfF�w�C�+
����D37��]�w�F�F0Z��UPT8�l��l@ݰKg��gT�C��OX��vT�E��VE9Is]D_���q���M�G��vi�Ie�����ՆS1കz&7J����2�����Ɖ�}lWw����ڽ��bEKĚǃ5V*6��Y7T#,k r¢M2�bف��	�r��0�y���^QD���D l�s�g3T��D�Q:]�%��iY��0%v!���o����?�1��s��39�MQ2T�~��Y�)�G&s�9��s���4��ڈ�ߞ�����af7�����;�.wHI� 1_����j��d'a��U݊V�A@��P��t��$(��2�{l낖��2��!Q!]P��`��\8��9ш%p6(��RK�֎�pUD�L����	Za)_��2�|q������"q��X�$ @�*0�^0��L�}ZL�	��"�`��P��Y�k���ā��NL�+۵��j/�L����.!�x���0l�i�E�{ec��{�]��v�)pCSpo5ԉ�Q��&�H˯�f'�n�i��]x��`XD�[Q}�8�M;,par�N��_as`T��>�E���c��{��3�Υ��9T�X8���}�լ2غ\М�٫D����6YGU,Tb�%���$���ֺWTz�J�Ael�͎B���ts�{
�.9{
sʜ���{EU�".����T̞:P΃MS�ɓ�xy�O�9��y���ŭ|�U�m�}El�j�\ϝ��k�������~{�KC�Ͷ�"���b"1��έV�������&L�9�^y��^lEw��^ȧ*�<�{<�{"'�Z����[ �g{ g�8���sh"^U�#(������K���w�+7����]�t]܇��uh)�"��ӑ�T!BY�0[J��p�Z�	ÝX�~{��=��:I���s��B�2A:��Ns�`�05���� T��Z���ӐuTc�Sqq��+ *"�*�7�m3���ۏ�OV��Bs�B{�����׫��t`�����1�-hhu���/oU6V�� Y��(��b��Y4�'�ş}C��|���sa[�k�Q��?V�j"2���%<���$���1?R�5^OR\��L�p(	��n }�����}�s�&`I�C�khK"�:�����T$�4�ŭ�&ע#�P������e����7軰v��D��=Ф�}B��R��:3 ��!C�ۮ��}L����1V� ��" �`29���J |3�+��6L@~��n�Kb�"X���yyA<�������w�~��qmf"bQ(=@������q��&L�3T" �O������=���s���7G:9�bq�0�v;�Ͼ>C�ұ0[�I��ə�=���C3��0g*���<�jҔ��	Iy������n���b�S	ˁԽ Y�#�[��
,�m�p����5������B"��%o�[�{��V���8�A<foKi��1$�eI��7�n�q��MwU,K��صz˵Y��Dn`�{t�e�r����En^o��'r�TO*$*�0���E���07��"�;W@�2z���ct�����~��3:�䣠h�v�Ά�H������'*��<��zcc2
� ��Y>���1Ȟ=C��a�z����f��}�./���pa���#���)�{�s���u�=z�=
�w�GJa/��>��"}���q.x�f��4��w�{6vT!A=�J�����%	��\1r��i�T����E���O�v/��<���9���@Yba����'&������	�>��>�������39�f�s��	���~{�~�K����3�:9�LV��M��#��>��D>a�N����Bk�����I�u����yh}�D���g;���Z���pNA	>�V�T�����5!6GP(g�|��yP�U��N�٨(�]�^�T�����׃��b��y������ӱ�<j��TMf'�0�I4���:\-�O[o0yYD`�t��]��j�=���cj�z�M��Wf;+�6�C���֮L�s�u�i͝+_f�̭��1v��_ar*Y�*�[IڽgV�ک�լ�$�w�ȇ������{=5�X�^�����O�j�1��BBA��-�U�<K�X��$ȉC�t��%��:��R�4<�\�s�C�x�>���q�`����K�,z��3f���h�j�6`˄��Ƚ�^8�V�N��*&�9J��2m�s��d�� zl�5Rr#ۤި�_�`=����`o턞�}�bW9έ��Md��������k����$�ƺ8s�9��84Dz��;�v4l��ܘi��t�!���%B╉HT�Y�r'���R���턆������&��d<$�#}�w*&��>K,��)����@;O�edAQ!cە�[>LuN�����h:�j�!J&{.D6�M]TD���P�4*������:�j�2%JOAJdc ���� �����07��Q��"ԗr�LҢw��b�B���yihKdLZ)�'P!� �:�Sǐ�1��I2@�.ޅ@��F��A!|
	�])g����$���x� �H���h_��;q#65�ٕ.�=��,T⢷�*�'wqz��6���;���׵��m�u�euꮝ��|�O2�s}���_,nc���&r>6`��-�����]�rg�ЈbH�{Da�#�Q�so���*��&�7>�!��3&Hh���؞�O�K?��?�R!��L��8I��	>���}O~���3��s�̙3�4�t�أO���{�$	`�$���(ꄂ{�+���I���v�����rn.�
%-�.��2	�N����.�V;���ψ;�XD�Ʃ^O�/����!B��A��N�w�!p R��׀��@�Y�ĆBV�T)��_�I�dj�\{����n�P�T)Q<`�9 J%�	�5 [4��2!��ZԢyl���	1-s��_O�:PA���E3�_���2���&sbO?9"y�̙2��l�ZCIEU�kGx�n���!c6�"(��]~剘�d"��)D�l��O,�	�62�e�{�}7\*#j�|2!��Ȑ$�a�s��`���̶����ų�%~D���߳��kp%�3>�1v=���E��y�����T&b��h[��Ǫ8�V�Bѻ ��y����g2ٶ���T��lu's1�c[x:�➧S�Fؓ/g�F�C���������T6�#��ҾMi���Ǹb�(�xD�<�g��l_	�h��=�:��-�E������Qg[m�7��¦{�);��O_Mh��C���QY�9^}g�{�޶�GV�V���<'��kK��N�Z�-�m����ww5�m�G���u=�yQ���O[�:���Dhɪ4^|����U��a�ZB�-���<z�k.;H�=�C֓�9�ɪ�k���q��<x�;'Q�Y����A�dl
�c�MKO'�C��gkm&�����͂wA�����<z[=��ê5� =�5��n�{ޣbDE� ��ǭ����-+K����=�=�=�ZS�<s�Ѣ��M6��y�xG���S��.�D��,�C�v�J�wc%'ulV1Uq�-\�TV
�����*,}�(��$�H-��\J"F�9�݁96�{L�ţ��{��h4^zi���G�����=_>�k,�A����1F0���������xc��������7�l3çh�E-d=mz�yy#R�e��<M�ڨ.	%��*5>~|��/�>6=b�l�_��3ƒ�,͕*��Ub�q6�KV����`�FR��
�{mv�F>�b�xɶ��[���҃�i��=���T=[Ώi��:.m����$h�n�͠P�4/,���_wDA��Kn���wn=������q�.l>�2�����!۽�a���M14�,�������s"����G��E����$[n��wY�M��d�9�ss���-�C��;5Ύ�d�F���,ӓ�����x˘^LM���%l/��:���&��ۧg>�(b�ĸ�`��ڊV�^�Ys�}�nM�^�Y�����.?e���N�<	�{mX�Y�6��-k	\r�r��*kw��M���G0o�`_(���a�9��lg�-�".S#k#8Kj�yyW�'r��uV/�F"DbQ�N켪���5{f�ѵ���ES�:�be���++��9�{�DD{���p�TH�/l���h���tJ�G�Q8UUb���(4��i���ӥu^�=x"�� �9T]Q����3]r�i�6���6u�ڋ5f\6u^F����DMH�p����L�QaÞ���� �����+�U�\VեRl�R�Q��m��UDNm'��w��{�Jۙ���Q6֍&�m�HУh�D�^�&�Թo�΋KQ�H� �m�1nu��ڭn�M�0�h��J�X�+ngS�:�Db5��m�ݐF�qN8DD�gQTdW��J�5��-��+͊��Ѷ������+͍u`�^�"�z��!�G�9;�^���ڈ���L��h��D����TF*#hȎ��ˌe��U�Dl*ʙU]x����DE;���31z��sQ�Wd{�QW��T�ܸ�usg�W��sݔ4��-םm[]A.���)����i��EDww�R�B�L|����鉉��|�͂�t�yͷ �}�˚�&���ތ��.��ܼ��GiҮ��ꝡbr�Zr�/f���i��x����}L��^j���+W))��!L�e�\�u�۷�[)i�v�nVn��2�ZƬ�WF��#�[T�t��V��+�p�R��5��NB��t[D�>w�w!��g�j�]�[a0��V����Ι��)��Ը\{���&70U;��|��7��	sTۭ���e̦i3)m����v{�5r�*K��-vR6�V�1mq�iب�w�{Hb`���9=���#:_ya��"���f6aS7���3X�SXF���e�C����V��x7�}=�?�>w1�H��/�Td����V�d[�"2-� \u6������F�r�S*���ڱ�U�96�ȣj5jb�P��L��ک�[���P��0�!	!pj�˯�R��O�g��9�pU+��D�	�#"1cjgPz��mD���s��<�h�a�s���<�<�6�r�׹�����\!ԃM�쳰��9y'92Pl���)J��\dN�0�-uZ���4��nf^����yr�0��9�V*ε^�"��:�G1�ʽD�{�'��5��E�[ ��uj�u��s�xj�������J2Z���Y���k��[�;�s��7Y���z�]F�k;:��c[�D��� ��޿ن��F�33��3&J�D��j��I�G9�pQ��6���������I��>�1�1��B�U����6H�-�JXk���챆7@�&�����Ϸ~�w���!�=$H3��_b�TM~P�cT��q���G0�����'{`}0�4K������^�\7��}uDT��
r�dB�����r�z���;�G=��1���t�ڥ{�W��<:I'�280w�k��,�h}����VB)D���$��R;����8�ɾmjZD>���d�-�ٹ�CC�S�(��À��$A3"��:�qǲ'h�|U,��)*&�Q��ǲ�xuSWc������8��+Ț<��q����(FfP�d�a�K�I!���6[��z'a�RX���`�F��PLQ\��ؼ�f�@7���h`Uq"g��_z�;�D�`���Ե �^�0R��� �� @��_@�F �鿑>��!��3�9�s���6q��������(aطX-��3r�L0ʁ�:�8�v�Z��)��gb��Җe-Ke�]�}d�\;DƥA�>|0Yf0A�v�j�uk�u��bYwʾ�v�삺��"^r�!�"��4�v�}����*����*]�d�]�'jp�چ��Wy����5j�v*sf,���<�����o۝шZי��������g>�3>�e$.#r�yQ$5� _�پ�*�xvD,(r'Km�X�}�Dy���C\�/�(fϯX�hR'�7�y�{�ܨ;���)�P��沶j�3��^��sx��A��6�ue�2F�&�|`M��웍�T��<���ŕL�%gt����}����$�S9U��w�X	�#"�"s#2�
bx�KKK-�B����^f��z��忘��P�9����ߢ|��C�丛�ՙ1)r�P�עK��+pN�bx���l�\V+���3�i�u߿_(i�k���{��90��@8��?�Qt����
A@�(�������U��:�.�T�5>H���NgV�'X��8�^���}Q��А7
��d_}Y���6Zc09��LA�]|4R�>��'���K��SӘ�4z�\9�83��tdTF�a"TB�
����:�Z�N�k��L�o�Xa���a�G#�n��j!���A0�Rz.Ϩ�D���������9ou�LmM��w�Z�91�S�э/�����lC��5���V�m���H���\^]���yATDE�
��s�����H.���(����/�d3�"2B��򉆧�`�3�="/�w���k^�&�4RA��6鸵*b�	�5��nH7�,��Ӹ=�o�3��b�>���sPT�a<�I����D�E�5@�l\Tm!� �.�<��k~��{Z��	�O��T@�Kʡ�)��&k.�(���7���d߇��|��*5��O�B# P���E�ˈ�5}TS9�s�8ᳵ�����O����G��$�4���0|`;���@�d]�G �Wh<* @��B��x�Fu��w�ʀ;*���PN'�"?��l�Ȑ�a9J*��:j��������]dU��zy��Xnqb���j׳12?}c�Q%㉋ �S	��[���kD���e�28LpH�P��IKsI�����5�A�5�P�Ǫyά9uD�D��4��($(�K L����%��i��I)#J(�%*��p.g/c���n2�/��$���+ٔ��P�E�ebvґ+̈�a��gz�Rǚ*Ų��/M�V*ԫCĜ�T��d֣���\�蹫M��,���9w�6�i5U��SS�b� � ������{3�D9]P�b�>����h`� |k	�躀�t��Y�SI7:��tg^{P�vDe.���U�A.ɫ�\A�ެC&���P�c�<P�����69��p�<��A�?cA�d�(�
~�(��(�f�h�=7�{��1��֌���؆`��s@w1&h��}�1eD1�bAP���^vq��@uC��@���!�P[�9[0mV\4d�D٨'7Jfs�:�x68*'�3~���y�sѾV"��Ճ����@%R��*�13��bBb�6�����`n1�`)psR�G���TO-��������`�iA|�%��vr�}'q����tڮE�N�3�%�>�.E+uȎ�獟>,��$ �R��O0���ϣs{y��"���5�N�H4���}���V�}*�w���}�ε����%��R�a��6t0QE/�4�E�5�R���xs�	vMT<����6}��O���9ғ�$G]�I�X���`-��)D���2��i�j44��pT���a�D�cF6���j��D�9�uj�yi̙�7<��ӞD�929c��8���-�)]bû"t{���1��h�G�柟⩕٪[�B��y�0��|1n�f�(�kXy�|x���[7QoEK6Ua �ZPA����b�95<4��9�k��έ^V��U�Qyܙ�7/`�r�9b�d�����F�	�!�F�,��9�k���{,}z�ʹE$�#�ϐ"�)G@��������^�Vv�b'(��in�q��kY��]r�x�?P~A �D$D@>�;4Y�aA&93�93�j�H�P��ɀp��{��90�8�!�k�է%)-p�CD�B�>ʕ�Z����qfŠt?���:�����z�.�_?���})P`��A�� �<�sF۠���9F�q��`�꠺=HT���I�	X�+�g=�B�#����$�'(�l����`)!pq>H5��O�x�VqټĹ�!߫���l��̎��({����`Omj]	���4��=^�ǋu�Q8$D�CU֕Y�@{��U@�	�a�x�6BdU�����_D.��\�{x޶ē$���C�)K}I��V������[�DuD�cOo�Z�m@t0��ApPq��c��1� D����*A��)��Es�=�]��r���%��/���7�׆��.��\��-�0�Y78��鯍������ QD~�@�*/ӿ~��8b�ٙ��3��g&sNֈV1�V�ʄ��q�B��xP	Q�d-;X���I>�zf��"�7_a�@UeXB�M�e���Q�����yH�P�J�	�J!J��hq�:i#0Oii	�{ (����nv�ϫ����4Q���Y��������4<��kN+�Q���U�s*�y���^=�R�F��X�Ͱٴ��{{�� D@Uu|޻�|��ڬ|�5IJ�"zrp"vp�r�f�$��A��yެv�>��ʒ�l��B=$�"�H8�	̥A�H�kv'5[�K�D�kb�TFS��Q�\�	X�xnXU�LN@-��5��hx��L�0a/H<Ȑ�B*�5��ES�D:�ߟ9qۄQ�U�z �Q�@��$ZTG@S����RϮ��Wx�����ɔ��v&��:r��i�
`�l6�0}��hO�v�f��ա+��3C�yv����un~�yAdT/Y��� ��┝�	�&����z��K���LB�	l�(KC��Z�3��Ί��т	��46�ϖQ|a�'93��6q�#��o�i�1��	�������=37�Z�'7J:�S�6���ب��h-����z�D#X�PQ[��4� qD'� ���ΉP����R���7�~�^ �C�*�qRI��.�v&�64}��\�ɯ�AQ#�z3v5���"x4,�>�k��p~�4D��Cqquȵ(g .� �u�{�ߥ�j���ӣ� -��9���:���Nk���,������R��z�W�6k��m�,�>^�b�N��l�,�4I{�"$*
���
*��"9�yߺg��������t:���Sċ�1U�WT�����HBX-�fh���T�'f��Z��!�n�y3]��)B/w8�&���J�L!q�Mm�Nk�Z���,�����ZC	(pr� dݎ�٣1L�;��.�w �����Ϟ�@N�"$.*�Π�f�f�L��Z>��) T�辇 _��g�����2��yɜ�92CP�dF'��=�~	K��s0�gG's��9�Ɲ#�����$M�XY�u��$R�`����R�.J��u�Rx0%c4�W�\��|��������T�b$�w�}p<�¡��,�!
Q�@�)h>�3�����D虧��/W^L��j�"ywT��p�s$����gIW �h��	��k�ݒ\gW�Th��"���Y�L)Z�5�5R��a[�.���!���7.�ٖ�M2`�W9�hyМb3"J��"��g^Q/5P<�B1��YA$�
�J��x�����,E%��[�51���+֥��%=�`�Z�˸�ۍ���#5�Z�ex��=v��4�M�3�d�WR�4�r�S���6=�n��\���>�=ƗXk,�9|���"��	 *�}���n�^�����Ԏ�g��!��2��$A�s��f�l�}�&���B%�*'�.�7�r��f�$ * ��y}ډM�F�����C�=���� ��B���uZ���2f!F 0����<���>�QD&pfra�4;[�#��w�q����n�N�C}�O�^��m5@_�!/b-�� ��[�Lл�!����ͱ{^��u������A��L�xķ�H֕UUUA^���{�6�W�{�P�5�C���&kZ.v~� ��3��ZKBH5�����ܛ�ux���Z�]'>$4cy2d2loRr��]J�{U��R��LM�u���}�C�y�j� ����C�f�pC��IRX �(�L��RRGa(~�D�AsY����W�<Bv.e��Z�!P�2ˤ9,��(I��b�&Rj�����cy�� ���I�M���p<����`���TOP0��xZ�@��n�����47]o����jA�3��ȅ��@�\�M���������������k�FDC�D8J""���������51����MZ9{<����iC/d�rr�p��9u{�UmEYKIh�çe8N��8���=�Eg��E/oB��q�\L���s]����}���HA"0F&��ծs��T뗡�riEs�3�ɩj�V���X+�+�/eLޭ]'Z�9��l��L�3�D���9�Ԣ-���s��SU�EN�V���9�D��u� HO	�ٻ���4�;�Q��������w�k�=E�P@ſ���-Z�ÄɈ&{��X����&s�J8��s��4�Qa zzh�I(a�G!&GT@�3K�Ժؕ�O��ƪ�h�	ڨ:ҡk��T|�������@���gx�o۳a�!���L`�%�~�Й����R}���y�\�[�K�6�X�*C�(
�tV"]}�D%B�:�9�ǺP^�v��,�O��9˄R��L��F�G�D��r�a�6�|�y�7#�=��Ѽ[�ٮZ��X:*�r�Q�`[��A(�!������㺩��pFD�y�S8p�gO(� 2?��Z��>�{�R��C�k�L�#�x�e��2��<Cާ�3I��UM��w^��O�Q+Iq-��I�)��e7A�3�3�Y�-�"(�(��#�A���՟��8����9���p��<c�G����Y!Af��l�>z��~I�u<�c��\2�ꃀ0�ț�����6fn�Gv��V2J �#����Q�LJ�	6LA��NV����gŌɉŹ]i}�s
�=Z��-��U��w19�{����Z�Nfn�imO9��k���9���{;r� yP �eFA@zv�vq>�)�OA*#�-*)�J�(��?���3	4��#�wP�v��Rr8�P��A}�g�I�Ji�֠Sz�-n�Y�S��}ʥ�w��'}	�%�LՂ��`�8͊��t`i��I$�P0Z&�5��F�ʫLp��ѡ�pzȀ���ȶu�$�p%mF̻��Bq�*X��=ǎ��$�e
*�V%��&:{|�~�{���a7��KJ���Ff+]��^�K�5����@�Z��,AFa�SØg:�*R7����{��=��fL�3&rb%̔�P�a�����!D���p�����{g�W�ݜ��a�SȆl�(a9�TE@��|Ok��>��c���ِ~���ƌ�,��֓�L%4Ǒ@�g��Q߲�y�U"�G/�T�>���l�����T���!���h��8�H0S�B�Q-/�d�"��]�6ۥC'8:j��+N���o#%���U�Z#��T��ҙ�s�~�S��gE�s�qoہ�=����9��$��x2�vc(y�nd5*��̬�lMd�ũ��Vl媚�%{72�,�'΃�T�Ws��\�����|��;ٮ�C-��h�2K���{GqW�Q��wl���X����Ġ�6��5�J�j�de���R��E��,k<�Ƴ
�.�C�g{ٳ׊�ʹ�ˍ���vm[V�)U�������w[�/b~�B�T#��rhI�ہ�38����55�A��N3�g�o�̧Ҝ�2e�"�h��o�8�2�7e��'���C����'�ᙴ�x�Q{mkvZ��.�j�6�G؜��9k���315U}���S;��O&cU�֭��^3���޳SS=M�ffm�A�59*��j�nd�����=:-+Ϸ�r���3]Ur�ʫڝ�h\w�}���l�eۻ{Xu���w^c�N�g��H[�"��ϭ�r����]�g����[|Y�~�w1F�*���T��V>[��6ʱ��4��7��fd�U~4mf�ᮬ�p�ϓ����Q-k�k�2��\x��.4&Z����Tm2˽�=6Ŷ�W�+z�]N�)oT�c����n��t���l�Pc=
f�L��0�*E�2���CnE�4N6������;��2)�(H� \T$Y	ut�Y�{-�,j���c�S�5dG�W�R� �t��l�M�R�mՎ[5fޖg"LV�w6ܶ7!�^���K8��xD��з�����+Yr�ӊ��]����ݓ�c�}ϫ�=dQ�eez�)]Ps�1�>+#�%z�ių	��i����dK=ӂ!	���M�{˱�Z���j�
M�:.���!�8s����ۓ��;Xidxǧ�cg��2�o[��h^��ݙa"��n0�<�_5��q�6�wf�Mj��w7gw�e��&�(�D>�!��т ��{ʾ�I�^7�L�:�9�9�9��!V_?=]�0P�Ď@�������rᵼ�S^�R���T2R�]��J�ܷ�ȩ�#K󸇙��2�)�~r���ZY)$�1(̃ R{���9�by�73TU@R��n�P�����F�������O3��&Y�&��X�d��z�AHT�=�d���4�*2%s���r&�f�[��{�C�8{xx�^���}T^�vP<�X�J%3B�%^p��U����{��xC�J6���)L�l���X:#���4�[�.r+�Ѹ�ov�F�S��<׸i�w�R�c�#mf�w��L�dS�^�V�����k�|��D�+ٍ�.P��Y9��)���6h��\f�(.)����U�����I����y���$�ȑ�Q�f�d�63~>?g�E�y�rgG
��gk�c�[��9΃���\��xӎG�;�߼}>�'�N:p���T?v�:%E��,�Z�,%�$�7�o<"MR�f�=N�c�
���TD�c��2�H:z��A�k5�/�Ԫ��9�ͷ~VDA��Ǡy�{[�ݷ�ȓ��dĲ��K�k��Nw�@<q�9d@H-���͈21�tA�b��ث}��������J��nӮ���hv���
��㣐�#Q�`�_Y���ј��3�syGT�{�J�茴�DM���e|��+!�a�w��!a � Sʄ�%M��� ��ub`]�������C���7��
�q�q�Y����d?�<~d�@�<�.Ɗڶ�b#Q�D`�:����urj�@hV�0Ք^�9���f��{0Dz���砦]ʧQ��UDKG�����%t�����3�=�d6���_~��v���J��{��0͚�/Kxc��XX�!+�S�B�Ib1���Q0��9�fr'W���y�W��nre�UU`S�3��F��YNT�rs�w4�3��w6�m�Α��vq���9�=���9弼�����Q��� `��"m�!hI�~��8�y��I���&3%�&��[������@�XI�O���*�/��s��2T�SSWG9��3��g0ѹ��A+'�������������>���T1u�D�\�<U>�K8�&/r�/w�=-Ѯ��jH�a���'Z(�f	����w麡�?i����{�z޽4ѝ�.��g6l����%V���l�G|N�ڊYӜOr��x�&Y�-���Ṷ��}�ֻ���}Q�f��>�`;����>�z>Ά�:��aiq"��H�T��t�»��z�C=FK�����XR"����ʍ�=�zn�vs�b�_�HN��$a(��x��D)�%�̌q29g���UG���t[f"
�� Ⱦ3�N5�� �L:����ĕ���'�V!a�BâN�Tc鴖��9�ts��&p4�'�z�������t�B0�H�%J8n: A]�Eּjې�S����]�{3~����CUʱ1�q�ͧ��G�$�����a���b�4�����N��'p�/�3$���R�5���uG��y��d��ra��o1�j�Ș���2sv�JY��}����DG�"�e�Xn_y	������-�"{)Z��,�\��_?w��)c�����I(�([�9.Eh<�e�2#̃��{3�o�������� Nc��aO#Ӥ�o�� ��G�#9�x#�n��e�|�`�,;��c����P�n��M=��;׵ض�7��D�v$,��a� Q6�LW��������u�,;Mz���t�<fD�Zu���x̅RJ��7px1V!�Hxgg&p9�X��&������1���dɜ��9���:1��,�JHG�E-Q���]�',U���Y�*�З�׊���]���D�+��8����@NT���ZB���:��ӵ��ˡ�5�B{�4z��=�l,��w/UzU}��99d@�cu`�����9�#��P6or���q֟c]F{��}]���������k��ח�����v�ͥj�Z�SLͭ�)�*�u��*�5�	v�� �ȫ\�n����e�Q+D��(��q�I��zr;�8v��AGݶ임��ݼZ`w�Vz��;���	�Oe,F��4NA�r R:����'�ӎ85%G���V���<�"[�K\�B�{���XdX���u  ���ՆJ%�����ϛ���s�Aɜ�3�����D���~��X�X�� po<Y~ۈ�s�݊n�1�o_�]��$;�R�A�(�h�H$q6ے��k���+��p׬���#Jǥ�-Z{��Sysv�I~�i5y����@�I)!)&�&VV3B*�]i'�o�z��}��&�
�gT]�cdL�}KCN�I	IUT9�j7�4Gmz�B\6�W݈\�"u"c���� �E��qč��w�󱓵\��5�˽6�N�����Tq�/NB���0ٛ�y�.�m��w��ve�h�[Y�" �P��!����!�A���s�!�[Jڄ"f�9�\և��tΦ�"*�$u���ّ�������o��1���� D"���3� �A�����QD�@s��3�f�KX���|�|�QH01 �@B2����=[�����^��J5�+�\�V�_˗�=^���q�O�!��$L�I!#��
����#wWD�F�ETW:B2����t��h�1iw-ކ_-m��w(&i��$&�����"y[-om`k�e����@`^t'=b[��ҽ/��N@!���@��˟{}�w���4�P�/�e�k������!�چ|�K�4Уn%��ǐ���J2�z^����n�[ok�3sL�a�==�sH�̠/�������� R6̟|����?A"H�����Tb���Ak���M[��y�3�^0�r����R(�1P�S���v����0����#9�Q��à6'����J�Ҳ���0�ά=���F�N+7<���o���o��6�m���D1����\����5��&q�^j`s��9y9j�Nb��Z-�s�i�"�ګy���r9���r�Ã#�p�Ύ��@���s��X��G �(�16��C�{������;�c�Z�髯7Z�ˑ���'2� �8���]�H�9��"1�c%�g9�gs��9���GHH!ʈ�U%�P�#��<�_���������IƖD&\ i�%
����ס+����ܖY��@��]��!P{ٹ�d��J�B%1{�Iyu�!�d���[a��1��$~�A�PH�粧 �C��=�3+�z�
H �T�f�8��yVkQ���P�ܬ��{�{��k���0 �)Ո;�l"��-Ų�TŃ������$�R&E1D0Kk�DG�w<���Z�o=����N�{؉q�!��2VgG6R��ha!Q�s�j�J%��������z�D�vp̙�f43N4eDϿ�)q�G�" ;�hg�%�y�=�:"�ay	bv>l�>���+��l2��%%�0Ǝ�4�������:}��D+t�Zw7՘�.�L��,ۻ��;n�+��q����m9Mu�1��l�V���FR���c�s�+�� �N����[}�mE6�:#5j����$�r}¼E�~��!Ȕ�xM#%$�I���v��΃�{������=6tP���D�Q/-r
��jD�|y4y!! �TUB�n/vV�k��-&�����Kg*E������E#n�c'(,��@���;�q@�oS��و���!Oa�m�V���Hp���y|t�i|�Cnx��}���J�93�-��:ǦF}O����:�QE_E��)�sLӃ�N�������>��>�5�yr%���_��������[����i0���ѨL]������I%�TC�a�ʁ=�/X����v��Ȟ�l�$��V�H�G�yL��f6ww�<�i�*x����Bfd�#N	4�����6\�<�듉D�ڳ;5�[�i��o�^W�ؽ�i�ݧ�v����[�Ղ�\��Q�gc>D6ojG�=|�D�����d�ƥBA	A$�*�Y��=r�'w n�oJ�!
�P���+���KO�*�����Id	G �ek� ��T�[�Ƌ����Vw��i���̅>��O��+��<��9�3�Q�M����rgG9�s�ɜ���r!Ω��Xb�TȲH�`Ȝ&�gv�zCwD�0!e�E���gX���N���[��B&#�i� ��tw�����툾��t�K�\a=y��dM@]Yy]�eM���z`�8�A�-��k����w��P޸1�}��p͈!�MRa�«�Ny��LLbTXFG�jd��~�f���\OG�P6A��y�A�������;�Cc�Cݘ^��H��L&=��=н��<��e�W�Lln�6�>�����mo������M�d����Q'��a��
5*&E��1X=9^e�}��� ���Hs�� ��h�o5F��p�9Щ��d9�����#�Q��@��(��EhQ�E���<�sh�d��9p:އ�Be��(�|��(���S��/9\%72����h�����0Ǝ�l����]V�ǖ�j�0�I�PxR��p����bte�m�*�MZ���K,��qH�U��Zc����0�/��^�54f�"q^�ܿe��c`�,@�)
=��Ǹ�����{5���D�ͫ�ry�Vc#\C.[�#��q̄�������O8�4�y�mw�#�|?�m
�GP'W0��n��Ȅ_z�!�U���4�"��8��JU鰜""��#*�gQ��TmZ�PDQ�?o�o�cnucm3/l�<�r��+�r��a8B��mE�i�k���hV"ڊa�W��<siQp���lDG��4QT�V/$`��J�u�"�pʉ���2/g��⎻=D�4hm͌Ե���\+Ŕe,&ND��az���*v5-�:؎1�4�]9Vr��4zN�[[��eA-m��<Z�Ji���������N��m���3���f�K�*�-���A*ҽj���;+��i�y�yJ�;\��:�;��o3����4���b1Kx��d����mJ�NE^_o>�TZ#��f��y9w3܇Y-��F��mZ!��a�Պ8\�å�1j���/Q�U��Ģ�(�.�ñ)HR��:+�@"ڪ��X�
�c�{޾7�v���f��ٶ�i(��˺�U�\�px��;�$�\4�uU��:��6�����x`��[Q�PD��c�w��ǒ� ���m���"-^��uh�`�'1�c���ݟ,�����a���-%#�D�Ĺͻu�׬��M�x'��'��OD���1)�q:k���_=ܦ̗�ϟ��A&<��eaK�s5���ڼt8��Z;t�s�:o�@F���~��1�������<,Cv6H���x�˚��׼��U\�ܝ��G�}�}a�b��ŭ�evlս/X[�-�6\^̝.�
��飃�����zJ;�����x�WX�3V<����ܼ,٭4�Q��/�;���k���ם�d~~=�<^Sљ�Y�=��n�w9�d�$�	�rc�9~�l��)�!�#$�lk�^��sgm�^nwYF��&��ܺj�'��JŴ����)�fDh��vZ�Q�GTET@iDc\/3��r�.\4Co�q�N�$(�Z�Uf#m.�l8s�VR�qV��%^��XtL�yh轞���"1�<��ּ�A��QEL=ٚ�Wtlcb0��(� �1KQ�*"�uH��ڙ����T��G!��d*"dL.�.�0Fծ�#���+��V��F#u^g4̒6� DW�1#��$��Ԅ"��(��ܵ��{M�8f��������W�)ʼ�TÝQ�J����7%4Fj7<m[A��[y+j�\����v3֋Z�eM��Q�\�/��uA5���27�<얣�{�2��q�DDN;�DF1�ޣW���s�m֊c쫗V۪���\wNEy�DW=�-�U���Q��Z�Ů��u�nL�5���؝N�[�h"j��kJ̻Þ9��K[��Z4K��[9k��k^y^8��qY��kӱ�	I8�FKp�*Im��N[lV5�z/</dA�6�����W'<+��́% �|���BD�Z }=37������l�۪Vܷܧ�ri�26ɣ!�v����22U����k7oک�B�_p��eݨ�Y���j�7R�kf��*�k5��z6�kL231�����ͽ�����[����V��^3u�GƺW˷k��{�xw���W�\�5��[Zrj��vwY����6�%�j���fiś~+�k�S$ִ�˾���]���ՓN׺��,l�+&=,.�>�Z�c�[k�MŽ���f���{p�L�,�`�лܤ�1����fF��;p�L��q��h������L���+r���/ֶ3fs���SJ��h���5BB�FDƢ������Q��� �I �kuZ��<��;Ec�͹i�%I��R�� �A����5[jmFV��(ܘI$V����)ÌV,0ъ ؙՐH��0D`�$dL#��(���:�ŵ5�3�%^�NL9��TN����NF��<��ꪠ�V+�*53�9;������/3����������	F"1ҷg�p�\�p	ݲ�xr��ɜ��� �pEV���r��R#*��ɇ0�/b(�N�^6q�KZ�9×���/=2;�G��3���~��qUL^sm��t�8۷7so�l�Ef�k1�����-��tb��.N��ؤ0`ǎ:s+�΃��rh��3N0�*=_�����	c"X�	~|c� �_{.��tC��N����^�W�z�]�"Dv���At	��`I�D��MV��4��-�S ��|-��̱J-Q�>~c��j9L��JI����8�&�����5>��v��F�C�OGP[��2�f�(�BȂRH��`Þպ}�[.���H���Bm:osQ�,e؎���}[��v9��O 9 vhW�a5K�����Y}~�@�A��Ll�F�{���a�},����s��Q�����i���}�uEBQ�
!Q�8������N>	m�[�9���X��]�C�Y�ݕޘD��1hy��i�$b1d%!2�Ju���c�B���.\��nƓ�ݛ�+Y[2�W�K0�t�uFC��;OZ�s�ʳf��ͳ���%�5����ѷ3���&3�� � ���J��s�$�t1��m�"�e-��{��:b��(�%���K�asy.!��[�=��Z�3~�|�lp�H�܁^TD|�C;�q�Na)�DX��D.�+sLW�k�Q<�D����;��d_{}��j�yބC�`�ɩ�"r A2(�U2"7�M�Oc�wvONzm}��5��l�2�x2�Ǹd�,2�$,44#G8s�Ր���q���>/�~\���	�9�3�"TD�����TIKG�J���ޕ�}[�ls���	�p5<5����\����R���ٱM(���H%=!��������{��}`E��6�e������{p<�^��֢}m��ɉI<��ノ�&���ʰ�y����ނC��uiצ����WCU���z�W��4m��W軖�#�ޱlm�l��ƌǍ˩�(�}J�i3kY��mZ^1��f>�׷y�?>�~V��Bg�$�IB ��x-CD���;^�d�l�&:%�4�
 C���DJ�@��g�룐�D�OC!��rARF�]�Y9�&�Z�
.��s}~A{ޏUX0��>�����B�?�-Z�9̙���<m
1#O��?8���J�0�s�ɇ9ɚf�a��������q��%#��z��|�@m\�(�8��#.f]R�TO?\� �{�P�V"�BZ�d\�"��8I�dOO��E�J����X��5��r���[w��#������CM9�4�$�I%D~��yӄ\J��F�NW�W�־o�Iq�����C5Foq��B$��E�d3/!�����=��j�L߳��V�j��Am�z��-uWݖ�żVb޴\=�y���V'Sp��I�j"֚6�6ݧ6���W�k##]���܆x���?!�m��}�j�~34zuO�H)��P�C$"c�����{�f�)���9ܐ�Fe
�A*�މyzʹ$�aE��wW�fL��8qQ?���!N������7J��#�:aɒg���1����o�
x��DDO���%�~��A��;݅o!�Ns�ߙ�|��;/	��)f���$��(
:�v�ny�vv*c�e�C��z���H�%]|&[��v<�_GL	�J<p�A �'��u5h��.�>u�kj�g�&-�=�wi�z����,�`cA�n�zy��yxm��v�P�#��"6�˻� M{Px��52���\�2�O�JHJ4��")G��h�*	�_y�"��|$sr%x����W�A�е���Q�/�qO�P"�*DC�D`������1�jg9�5��m漼<B��92�4{�p�V-��VaNm��`�3U�1+�p�!�d{�<��耑������PY$��%u��ѥ�s#�"qo�#�gVy�0��U�����8��#�k�7��c��&t'\�9�S�r�*��+���X�U��Qz��l������{���	z��M��mZ�9ɓ/'<�"����9�\L&�#jd;�Q��;W5����[�m�]�ѻJ_��S����pU�s3�935C"hߗ�u�=��l��a�F�[N�1�1��f���[u�x(�D���{h����K�HP"Q�z��J�a���!%���ޜ�S�<9�"z�E��3љ�����ɼ_\� ����GZkV0�Ȏ�~�ƚ��ܑ,����#	�y�)c�F�iO	����aDt�*�[�':���9���p�UcD�٩��^U���s�["@:��1�ޝ�w��n"��em����IA�0�!���#��'��دp��|�w��@�DN���O�w����?e*�8p������~�����p����EQ}
�|��0�4͜=Q����'�|1��p���74E��!
�a��2�\�
�uy��l�앥�� ��rlH���0��BA O���ۤ&De�D���]{:2p�Ċ�k5ڝ�V���][y���{�n��A3���}sw��/N��*�b��^�^��J�uv�$=�]�����W�TB݆DU@��m��Pܚ�7pi��|��I��D�"U~���� EC�t�m��n�9=�Ht��QbXL#��(�G(�!8� �z�\�\v=2
���8��c���#T=��u�SF�k��D���Ӑ�� q{�"}���������hY�ɤF��rseU�X:w��	wӮpƞb����4MÓTDD�Ͼ��~����;<�^�;�s�8:$B�e�`�BAB#�V���Za͑;�e9��������^��Z��[�=Z&q�BAL�CP��2�Zs��B��v��e
�
����Zoh�^��~��{p��ta�� �M$��$M��r�n���8���}�{%g���T�k-yZ���y/�Z�,�s���|=��[k�n<6�f�U���:F�6E��El�D|{yS��)._����s�f�$�A)c(�.GK�+�O��@ChۢL�f��c�w�I�|��3��g���4����<"�v�t�!�D�vS1���9�!�y��|�鹸����	M^�{a�!P�a��s�&
�F?��߯߿oHa�Kl���fs��%3N3�apc�>ޭtѴm��X'pw�P!*��W �@^5�� C�N�s����{{ճ�[����!����9"IaJ��Q�v|b��y��#j= ����]î\���B���z���A�����*����b��f轇P�:wh��j��_z}�!ڪy���&V{*���G�A�)� �=mȓ�E{�2��oF�!{�|B
�T#�tc��v�������|��4Fi뚜�݃5�q��U�Һ�m������Ѧ��=����u�ۻ�����-�UTu�y�{���۔a�;�tB�k)�U�:�yAf��Hڎ��@1�G���B�g��}�����Z-#��9.C�튑o�����g��k��ɜ�&L�3Bq��FY]�����>zSӆFAЄ��"mz�[lLz}sևkH��Ȋ	q�o��L�	����Q���zFJH0�$�RF ���V<�Г�Yy���8�G���l�(�>��ۖx5��S����:�XH<�	$A��Z<J$����G����^��|C���(�T�pF�Z6��NGI#"D��z�;���5�8X@z�z��T#��>�zb)�&��ŕ�9`γ�#�Da�G �|��6T!˓�Z*}J�wM�Ff!�达%��Do�w�0�g�V���L"h���1DcjڃB��#8D�s�W���rh��g9��;�'<�U\�i����X�"-�҈�Y�d�E�j�rO����`2ӎ?��/��!�ݴG�#�.Y¥���t�!�Y����'����h�~Z��k�c&b���W�m���<�`�R��"ƫܪ���<웥b�Xr��j�xL�/W�;z�Q{�YDZ��jW/e�������
����434:�=
�N.�V�e��V�5�7���\����*�����
&$�(���3t�s��)��1-������s2�;���fa��:t��G)s[B� ��AL�S|��T�kT���c"3�vc~/��פ�e�{����2���/��-0���HBVCrt� T=xظ[��N{�̪C�&0��H*���Dח�v��œvw��wX|@ݖ����L:q�b��"��'8޿;U�q�+��5��
�D�\��sD����wo��/b��asC$���0����o���g-Z��7��p����x��i)�Q2,�<�`�H��E�`f����譚D���(9�y󱵣�L�S��>54�k�f��g8+�� ���߿;�-_D��(�B>_Efi�)ƉPG��~~c���t� �cPF��$6zۛ1+�^g�u׳/��MZ���@�d�Kd�rA����
�,f�@�뉨�*i��{��|�uԔz�S�oq�7F+]�w7�H���f�|y�͘6�"�[e�k�ԉ��ǎ�����5lͅ����ٙ�����QId��:yEI!�Mg�koz�u��`��>꿙[.��v��#����9�����2e�����"��m�S�.����!�w,0@WI�SS��z���[�1�S��N��a�5q�q�-�4h�0�~x�j��^U�8B"(n�=!w�&�U���k&�����ra�fn{��J"#���;~Ѵ����Tp(��#e%LQ�c��6�(��Y��L��|i�'���		������g��鞘�A6�D�Ep��q��BBA�G	��L7W��o~x����D*�W���yP5�=���s+�Y���D��ţ�Q$�L��]/���$����G�����R3=UK�K�����[P�OE��D���楫ܕ4�*eܪ��7/6o�^ⓞ���FlB�D}��ټ��l����V���]�z�X��Z5�|��̘���8r�gg�3�N����Ҷ\�L�[kvk�=̓�S(ϙׅF�8��3��^���Tͳ�5=b���eS�Q�{�����CԢ���ڝ�Q=��yv�wt˴�y��.�]JҘ�+[pK\9E�d��(��:�u���j-F��biV��\<�ջ������x�����s<}�����4��d+K;>�F��Wo�fںmA�k�wP�4����k���������4���Q��-<M�%T�ݐ��X��H�͙Wy��3T�{&��1j�����P�[�em26��n�uxTH�L�﷒��{�=6h����y�𙚔/�f�)>*�y�jԫ6>KQu��JCl);�[/��KO���T��l��5��
F,nK]��l��׫�o��j���6��d,Z��+.�7V��+qh�����yz�jk��|�h�YVlל��w�#v7uvw2�cIk�Yւ7#�֓mr�fu�׈}��]�(u�
�{e�l&[o�q�a�i���g_z}m���$��V�YWn�v�n(������a���)r���c#G��raMѦnJy5j�f��-��uV�k�h�Z�����˚�kY��r��r�
��"�ɲpc�dK�� ț�P]�gQNM����Q����=-X܍�1ݝFu6W�S��\zvkj��+_g/V[�� ����٧�ms33���4�~j����j���N>O�D��!�_*���҂�'od*=�*�2����Y|eDUU�&x�;p�R�pr�% mzsQ"۷��y��C!��B����;�@��RM$�U�fXx�QE���An��&QO�p9�ݐ�gL�8�NG�����D*�9@���h�<����ڝ�`��q��i&�b=����
Q�Ҟ<jP�A ����ݤO{�.��m٦k�thAP��>��`��D���8LV���Wgo�G�b	$���n�%�v1Px�����z6vV�"}=���4GX�X��Iy�Dj���b�=S��:U�AF����DwJ�溅:����v�37`��w�{>��W*��U�|�3v��[b�v�fgq՚�]��s's-e)�3_#>ۭ��;��~SR�(�� gCj���'="[(:ۊ����"[�^�&�-��=�	�fT�x�����f�2g�!�h -رS�?�a�L} (��L�4�4�D*#��������A!
&6�4w�TS�$d[�Ȗ�VX���v���_	�J��f@VʃL4�!$������@����z+����qL�7��-�K{��2C��:��C{�!'0�:(�s!������Ym@,R�{5Y;"f��y<���F�'���7��hEBLe!	�Q!� j�w!�rM� �pesH��q�OSVd�.s�� ��,9C�9�
���Ч<Wz��u֜�נ<K��Fc�����?�!�d�N�9�mm`��A�8e��j2[hՌ�TF#FL9��������򝞽����NN�ѭ]�j=�*")J�J�h��N�za��Exc�8r��1��4�e�Ƚ�ǌ~݃��kZZe���k�ԙ�! Aa �-�S9�m�/drj�{���i���+�!ܪ*�f�3�f)�w*��p�9�9��8s���-(�\�fL�x�s�	�Qy�r@��G�[��|ϻ��zoz���ki�e颲�u��n�F��Z�{���O�-k���Û��+#�E��ɣ��i�r9�6ki��#5wڿ��=)��^ ����e�y���H�N�F�@����!ж�af�՞ٟHa�g�~�&ٺ��� PBA��BUO�/�c����z�Oz�ª%7<��N`TzcB"3ψ�����o�$-�A' Q$�$H�(�D�ӓ�o4m0����5U���������w�T�wt��L5
*  ��=!Q9k�eze��н�=�<Ҧ����y��ű���/=:%o�u	W<�ц1�� N��S �H?z_fx�^Z+�=A�Z�wx '4̞|>I���������f��׬s�g! �;��?c����(�
(�ɞ�ӡ��x� ��������X�,BD��~�@A!T%��ԍ�dB�)��������vƕU�'W����dɐșIQ%g�V�����,{'u����Em�\�-�+�O=�4N-�ˑ8��Nc���1��W���Nܽa�[+Y��_��n>y�w� ����;��}�5���R�����ZqI(�:H��hNKE��`�5I낡���s�s+%ؖ*���/u��0���7�M�D{�j|���0d�w�dO1��@N� ���A=�0�m�.�n��O��p� ���%	IBN�`/�?p9�g�Q,��ƇG*��y��D��F<�'�2�}�k�A��b�Øh��4LTȘ�/S���A�p��s3�&���CTA������[��"چ���'?��B�<�\�!5�����x��Ay6�k΅�%�A�%�����Z;�X������-ۈ����h:��.�.{�����c2�v����H8q�ĂA�y�Q�`T�b�X���}�'|������1�*�����6چm]Ѧ�ݲ�ڷ<@�Ďѹ��һP�
�X�C�����.�Z�J�?y���tc�}��,���]0�|jjT�A2(2�_��q��߱~����t����o��a��>���a�/Q5�[f�p�� ����	KhXèW�Ʒ���qx`n�D�"j��C��DG���0��k�L� ]^�;j� 	��n�����|��E>!GS!��Ɏ8D��o���~��"a���8#� ��,���ֳ���Ů�ʌ7�� �!�3r�!�FEX1
�Fs�Һ߻�v��=�
�M��lՔ6��C�!�a����S��Bqic���* ��R'���/�&r����!N�x�W�����D�8EW<t ���4�d�pZYB�<�w�����:ᇝ�Ca��jf��{Є��nԾ�دKUV��3��R�6c�BSz�v�7od�\��k�|��2|4W�>�e�a��׹u�����
�1�V�Ŷ�u���5���?�;!�
0Iqψ$�x.�cP����2�j}�yvfX��:˸��5SF~��
������o �}���N�0(�� Q|Zhaϒ#�0��$7~̓ � ��&V<�5<`�K��Kpk��ڽ������qҫ��A���N\���JI)2*��#�ㄜ!(O�|Ǽ��k�P���
��B�֡()T��eu^�e�"������s�i�C��*kcCV]j���j�W}��f��˪B�	SXؼ�bS��d��H!�Cq��f"�tG��>Y�����S6�(��|lk���<l�r'U�-hi��I$�G7h&lyqY�#���]�/�R��?��\{̨Z�|�wu!aCX4v5k��KH%-R�&�L"b" ����:����F4�
��+4ffr'f�<9�zًr���n��쪢-�ݱE+����<��8���(5�y�iQp�zf��2<�u-D����N�k:�F9��u������8n20����j&F�!��8S�r�y�]ܼg�ʨ����ީS=��ztj��<�)���x�-j�C�Ƀjgt{d�Hr�s����H�.F�0E���|)č9����ٲ��w��%�������$ăqHFX��hh	�:�F`fƤs�����s��4�N02TA�o�?���D<2"9	��]C� U'����
�7=�v��{��W7~Cxo �	ُK�qE�A	d��"!���9t��_e=�M�, w*h^C�(���D�پxǹ����k�x���KB	7��@=��9�G��[m2�U{")��=r&�K(�'��I�� �B�K��mϭ���&3Ѩ�'�X�T�l֤�AXh��ghU�ӾN��j�k�]��!A��q$B3�z�<��Z�3G����7��o,��	WD�{�v��D�ȏ����<Z�A Ü�ɳ��PF1��������Ѯ��G��gɞbq�W��߾'>1h:$��y� ᜾kП]�t��������g������1�'�pq�*�ƪ�Q-V|��S�[�o�ib���R�-J�����M��SC��u֭���U�^�1���k�u+N��>������7�ӱ�W�ZѪ�K��V������~Z�'�)�d:�+:�̭7U�x��*x�R� ���	d�(�����9 j��{ٶ�/UF&�`'%�P�!�+�ݻF�L@�d�T(�����>�wE��d	ETE��[Ӄ!��76*���Fk�z�X�q�#�21C�#��'�_���yv�����[��D"6L�,{X�DÒ���QB!�`q5
0@��|>�A�������������8��g����8������-(��� ����N�sP{0G���s!�$v��z/b�ge�![��^2'I�p�zID�eUD֡�&Pدv���L�H�,gr�"e\�(F�W�X���=95%�)c��砊�:oחa%p>WGNס:�5�uW�����L��2��fL�"����]\\Ľ3��^�*��W��I���q����7���q�^��/�Y�dT��O���_��#Z�X��4Ddq�(t�>�J���o���:�]�n��d=WX�{}��P�:e�W�6.�rI$��&@m���A<��f�h�_��P�u����J�FP6vܐiȰ�
D,#CB0���TȚ~��}�����wl�ɜ�9�i8���'�����RB�! ���6׬/���B�-�;8B�ɡc[����G�+�h�z'ɥ!�&! �H�&��G�J�ov���ޣ�۾�}��ďi���V]b'M��0sF,rA�@,Uu_!���G��r�|��syP͡:�	��j,�C�`�x<Ȕ�˯������҄��g���E��Ef׎��z%爯K>�`�L��Z��0�W9[�t���uP���_m�FYƼ�;"�FV�R�n+b���D�u�{v���M��i	� }	�3sA����d�[Oq�	��D�jC����j#{(�hL���?�XXb���3��ڌDDo����F�+93�.�;9Þ	0�A,3b�W�� a���<��8N���k �c�	��*��6Ŗ�|��@/@E��h�ᑉqa��/3��$Θ�J�>߼����z\AQWHoz�}hwN�I������	�I	�A)((ꄦ���F����=�?6!�['�g���5Е����K��;Ic��8�#��fy�)�����L����U�{CT/�NZ��N$�{~فb�:��F��k�@ഷԄ�.@�@Nl�`IS�C*۷���e��`��"�U�u�d��(0�y눈��t8Alj�W�6��*0˄]Dx�U��tx��2'6TΣ�ũ\�նˢ/g��0v�:�&�4z<"g�=��q��f�j.:c��Ƥ��iF�����QKX"1]��"�w-\r��z��[Q�������5F2ƗV�L�4D�s\�����J�5do'd�DF؏5��X�c�=�D�m�X�,��j<',W���.��E�z�%�T푭
klA5��Z�UV.�{af�4y5��M\5����9��KGT�� �(�ꛫb��9w)��gF��Y�Z6�k���Vܛf\jڶ�36�����`qF'#Uh��=�2���ˁ�����2���p$d��DAE�^���A��sҏS�2�^Whdy�b�Ub*������� �mETUX�66���v��*g�A�gX��3�]��Q�Nj����ݻ�TWD���k�n]ɁKc�5�-FD5�͋��؋h�-s�j�Ճ����*�M��F$��Mm ƕ2������mj�3���W�,v3��r̴��u�2��*ӭP=��NC�YyiN��Q�6���5ك�]SF+�52����o�U���e�t��͸��|0���^cӟ�z\9�D�7���+=�آ�����k��qb���n}휉��ϖ!�o$_p���Y�٭fj�/�|�K1�١�'Y�݇y\Z�]��%��[�k����i�Vǖ7gYYs,gy�����2e&)�zWn[ZU���V.�3�Z�Qr�k0'mbr�Zb奣jF�m)�fo�Ȗ���ո���بej؊R�"�p��h���X���ic]�d����"^՛w��''�N@�{�v��ҍ�g�k��nx�V�[����	��I$����v����9^j�"B�s�y���eUePDUDDi`��cEf�UG�oa�c��b�*�^�(�����*�y;��Ղ"""+�X�޶�h5�
����y^��*���DXU)D�Eʫ�\��j���ν��Rf�UmDD�W�c��m��[ڪkn�um�jՆEܽ�mZ�DͶҶ���6��Qntsg�I$�d�50�#��1�"-F�m�F\�S��VkDAU�#�j��x\4��GTF#�iVьFWQ�jdΣ*.۠�#-�k�V1�����evy�F"1\�7��X"��t�z�DDJ�ήʽ�Z7)�����ѥD���W����W���+5�W�lQT��+�*HƸU�g:������ �٫P5��x���W=�=ͧ�{��.yɊ�*����������ʽ���ڥ�V��)ד���5�ɘ�.{�A�ڹ�r�QvH�i/<��ޕUD�@ܑ� Q&���	�ڟ8��C�y2�*�û��Q�"�;5�5Ow�:��Z�n�s���Kv��K��Wqz�{M�e�C4�Nf6���s:�NU/e5Զ���4�JN��-�;��ͺ�[5��z��bKc����Sj�E��s��r��m��-�l��ǻ�?��sU-�bOݷ!�F������n{�����}�S��D���t��S/���J�-�y;0ӹy���7��,�5�M��nV`��Q�ҳ4f4dn<CKe�dQ��D��B�X��O�s;[x�>�;+Od�*���Ȳ�p�`�[��W�q�N�|��sݛ�)T�!�J>�?">�SpN�S��DqL̑T*T\�@w
��F��sQ .(�5�jͺ��m�c;��6������E:қ��Y��D��i�FA�
ZQr0�F,��Q��V#���-�39ɜ��C"vy�4R&N����<�r����v��T�9y㞊p�Y���2�Y�z��"#" �DD�\��t("&���L�s�f�9�s��W.���b+g&fp���TUY�{��<���mk��`�9�nw�^aȗ�)�� �Ƞ�H�Qbm>���&fj�Tϥv]�w.f�hg�̩|�]�k|��_� ϡ����gݣ���3QI��T����0Ù�3;�a�a�WVBtr:�f�ܐc
q��)��"�ΥMJ
��s�._�[��y�we^�-[x��CG��"Q�٢��B�o�c#)��!���n����:ڧ��;+�Ν�˹Ȅ��6�rZ;�D���ǺB�=���f��Sw?E��\��P�D\6^ �D�]zq:�8 x`d������y�e}m�-�x��1�y���^lz��n1�]�\!�����͉�yED�" ��c�$�V�LKd�>�`V��ty�}��;"��Ĺ�2�1���ˎ����5[�gh9��A1"����8����&���8s�d�H��	�����}
}?�B��H�H�����!����;�_���f���L^�dǹ�T:i���bGqД�:@K̤EEp�E�nkH��7�=���5�C��ٲ�iK��~Rd��S�6��'�f�[/.wq�\]��ѝ�76q�Ɉ����Z�D�_��n��n�@�A���z+r�94a��&�������ܩq��#�|������������9,�oUǎ<A	8�d�y.���˹��s���1����Ή��½�����P\9���RL��Rڞf�ɡ�f˯M��W\�$�j��<��H�^��%���������s�8���""������6|<K�b�(������N�8`����~~|�C�0x���v�<��$�%��w���R�ne+��s9�XC�@�!�cMp����gy}�����&6D�vȋ:��>V�/��5�䮖ƙ�����Qe���B
��u��`xH@�e=Ldp�߰I<\�FD��X�]�\e��Q�;���y��ro=��LCK$N��&��v��s1��͇g�ұ-�k5�E}�e�[��ɓ�BZ_�F[&=�X�3GŤ���_��Y��Rc�jW|�յ�ֈ��/6%�qrb+}҇<����{� �E8�$�Ҡu�]�#"�o2�g�}�"����$���z��D]y�/�߇���$H��ςk�>Q8X!@�0A�n�n�t��(��ER:g�0<i����}��|=>��9�&؛^�hP�CZ*��j�H��w;x��{�x!T5)8��  ��>�_܁��~Vۺ��6���d�ˎ	|�ON@�0�n�R���d<J@`�9�L�N�kݸ��H��
e�5���W��Е�=yU%E0�u�9f����@ct�GKÙ�ݑ� �f�
�L"$P�"+tU߳"�-ݽ]�54T�;D��ysw�[�����ݣƾ7SY\�լ��c-C�52�:��^��5��q�lJ����	���K"�&PY	"���F(o���#%����(sW0W��q��"/T�߿�ӿJ�D�C9ɜ�̌�/������������L��$,�DX��߿�~�>�|6bq��$�}���x0=Z�1W��8^��Um�7W�Z�ܻł���]��(��Dzs��8#��[�ΏN+O�6ß��q|٪%m��,�5�5�l�Dq�a�A�K����;Ǒ7���� fhD6gZ_�-�4��O:�\��Psf�����a$�A��'��A������hf�#�XD��mr��<�파���CA�R�Q@��F�\<��~��{�}�2����|�B�-�a�&��Y�����0��95DF �Db"0`�9��k�X0��%��-�KF��0mp�u�^��r`i�iΝ�\�r�^Nd��S"��Y��R�#H�t��4ڣRgH�����8�� �?y���!���{�B��k��k�5kF6-�V�۵i�R��4��A$
�A
B�Dlr�CVƛ3������g9�r�h����j(���$�9"�!QE t�s�8WH��鵣j�Ç9���������U�x$�8�Q(�
C��22�h=�ӭg/�o6Vq���˵��j�χ�!	-��Rd��3��]X�"3��y�s���Ӈ��49�p �R���OD�a�"�j���斔=@z�'���Br��aZ�؈����~��#�PjJ ��R���=m�x!���9�����n�9�$��-���^D�M!
@��PU�|A�Y�2}V�\�.��VL�{:��:۞�*��L���Hq� �l�!��m��]N�j&m�QY8�.]d6����ͬ�t�.R�#U>{D���	��!㭁���=�V�W9]��-ڼ�ˢw�d�XX�ج�O�T�V!�!������TDD�z���z|�&L�9�r�M#2d��p�}��n�(��&���š/3��Ϲ��*��t�u�w2��]t����"���U��G��8�:D���闽���7"|����áƗ{y��g�j��vª&���mV�����3jw'�o���ws^%�$u��&�h���ݝ�6�]�"�g�����wo(�g�O f5@�y���fW���9���8�z�
CKDL�@��5�U����"��P��5S��9S����!�김��d��) ����^Uc�4�{��P�%���:U�[z��"j���/�w�լ�<�ȅ6�rq@�A�O���)�'�!-�ތ����[�����7?����ZH`s�7�C�����fp�uL��FЎk���6�hj�&#J(�QQB�����=s;~cD� � $����w8Hڡb��M�򩝳׳U�Y�@T�k��(��w� ������l׽��l��k�.��D�ˉy{B���Ej�����I��E NNr�Q�D��q<��{GD����=/�M��R��/d����D��\��*c^h�}���ܥ�ݥ�����k3woK�[��f7pQ��4z����s�~i~r<�}2��f��ZrrI$�D	�����gޡ�\�Al��H�A/�!"� ̖��"#6s}��V<���,�q�7���}��FyZ�������>��� �`-&�ߛ���ޔ*�&p���y�`�'K>��d�����(�Q8چ���ё�! h]n��"H`�8��A2(J�ڂvx�Dl�((����F�olt�R�ؓ��S{���X��b�9�A�TEX���DH@��v�vUl�C׷)|䩸���P�5[�s��{���P�)�d����|�ϐ�G7ف��L��m�le�������
!	ء&[S�B.g=���r��\^mf
��י��<��{��ɕ���1�oKE��ai�}3����Z�km���mF�C�ݭ��63>tnlv���F�/��mj�+8�m�����t������_�S�3J��H����8����9!8�nF���Y�9����/�|�Ot�Hh���ý4$�o� S;��dɥKDDA��o��>���&s����9Ѓ@ã:A��P()jU����D-���i�dzA�DF���9=�~����osF,�hiHQ!	2)J&�\8l��"�s��9���%�=l׬���S��-��b�LWKk�I��v[�32���v��煉��J�_�9���׷+�A���}ҡcͺq��Ѐ�=b,2����;=�`�'8O@�8c�^�L�DdL�[5oV���� �! �VA �z�����P����2S�{��W`����Y�=(��Y��A�����hhj-uD*aX�тJ4,GT��f��"�#��y��yy�	��&m�x^y���+Jǆ���N酪D�V4{��Ñ:�$�Ϙ��'�Aqo�;�x��[�q.8ӕ��vb��e��ffwZ[+��V�gvnh�	A
�B�
�A�$E�+��lkZ�-�헳�L�9�9s�����*���������cr'g���4i[x�uoe�d�жʈ�aZ�8s�9y����^�]�5�L�\�c�����cK���ǭ�ƼQ�Z�Ut��|�����Y���Ť�8VbF��&L���0�������M�;����ɜ9�f��u>=����d�=!B*:�?~~�g�xy^�#z"�:����oo��lF(���HS�f���Ј��j6��O��6��U{{h�U�F�׶�.���B
���A��������K��`9��X}��z��e�Ez�-�B��" ��B#^��9y�e��\�z�7��%�G|ʼ�ݝ^`�Ź>6d���D�����ډ��������D��$2N��Cٹ^�Q�9+�E�Xb!��x�� �*���7B!�@9܀q�s��c�щ�o����}��0X\BY$4����Z;�b�˄�|#B���}��[�y��̅��7p���4��0�HT9h�U��<�ص+l�ѰMU/�oQR�S�<�V�n�$(�]�OFwsqWX�j��ed��KTM�f��U�K��A��af�o�&X=�&��V=;�}����$�*dYA�)��$cV8��}���]���:v�˗n���M��F�O1��/+�Z::8�$��_g��'#��Q�y�	�D��j�E���#yW*��|�j�#Mr�郆%��A)e��>���N�t�^���� �g�C+ܨ����ɚ��tF�Q�0U HEe�@hd!��P� ����lL1
]��s���ř�d{1���0o#��((ݓ:;��oBE���g!����{}�9�{��������Ǝ8��O����^�E�ȧ��!�B{c��\�=b%4�Fcj��?E�Òr@�H!*Q�OZ�q3�[1[��.�:�AM�)���b���3�b���B��q��sww�D��N焊%��1��E�$[��A/.�.L4e������SQ/��*o9�ޟM�#/W��3/����K7��V��#l\���|�yiGۗ�[J������|mo��w�羍����d�R��}�on��$�c�D��{��+jf7"�b!��u�W5��z,�El{�yl]�WjE��*�f���j_3iel�N�<yČ��6_J�Da9eY����B8���Q���8żt�¾"���Q�m��5�:˄/v�.���mq�:�J��9t���]ʍ��*�ƪZ5�sr�a�Պ��և����SpW�foV��ra�ks7v"j��Zw_]���.j����!�]��b�i���z��ݍVs-dz\�w��W���|�ˉ��̊\������{�e�jX��مxȂP���Oz����X]��m�{�-q�Uy��,��l�j������5������v��tH�G�p�O{�d�GJo=-���c^����~+I�e��cJ.����.c]�l���aL������5��Tn�T�k���T���l��j�-S�8I��ɯm�w�J����������b�:��>)Vі����n�ى�gԗ�U�p���/�-�uwO�����A�6�N�M������$ʇ��VAO��rEvD�G31�5q~�����ő�7�1�+�ڱ@���L+gw,ܵr��g&�Y����eX�XrأQ@�Id@*%E}�8�{��kٔ��3Uk��י�����lʻ�}���K~�ͅ���DF&T�D}[��φ,�����@Qb�^�m�T�:'kC��p#���B��G�g�����+H��� s�U�r:������\C֮ٷ�{/u��\�"P��qhlv,�>�,���uMF5�ffs��*a��iKv��3�8{gp��4�84uE��?�����dH �@�^��z�i|d�'���z�
�XX�S�ޖ^$ց+���W�NOABI$$�p{B��Gt��������W��jr@�v^���`CL���Mǫ�'�HB��	Ht
4A�"i�Q1kh�i���%��1�ז��7������8c3)�˓8b����v���C����eZS؃'J't=�y�z2����D(�ѝ�W7)�j�T�\���V�i�ǵ��m̽��sk�V3�s+��mYsI�Ki�mw-�66f+�]Ջ�s����Q"���Ca�0upS�N{���b{���׶{��V؇�n�;ZB�!�jt�����$@�*�(�"�����3
�ά���}���V9���Q�p9������8�Ћ����,spJH"�
�F�3��C �k��P�?����^�{�'��H���c�9 ���������|7����m�A�o��)B#P��&/{�S�`�H ��1����C��,�.��%j���

�Һ��.�G!�PĒ�$$��(U!D���i����nP���2]��hn��l�s�gFe�`�o��ԡ*x��N �/�����)"P/��j�<n\�t{9.@�D7vl�M�_���R������	�䚭uDFA4D�D`��`ڶ�M�8F5�g9ձy'-�,;	�L��oe9�ij�nt���ETDH�eHb���{�z/<��N�������&y�n��p̱j�/z�Ց��Mu��}��9���c�� �L@$&D���3�ڵί� ��3��ȹ��ޫ���, H!NFP�%�I�7$������;q��� ,AIY�VԮA싔Y�C"�拙F�[��3;g���޼�6,\ٍxfwh|�]�gk6�V��r�����3����6��yݜ�p�4���?�;���4s�9��2<S38S�t0M8Da?������L$�1�X)����hB�;;��6U	lX��cy[�v~&c��Q/,9L��H��I)J)���@�x�Z	TG)��m�����K!�L�Mf�*'����z/qk}�!�c�A#��P��"��tD�����n����]ʔ+ޠ�Yי��K�r:�ލ.n��9���-�P|ۏ�%���	�؋�v^]<p��O;oEg$��"p��#��w��Ӕ�tTGs�x��TB����I�"\�a%�D��+�=??��겹���rj�f'LΚ7H�o���B|�}���N4������|��q�������0��4�	��TU��Ĕk���ވ�[Nxn��@y,0I�� ��I�|=��y�����=t��ٗM�G�_	����l�ەyݞ,ə�1�Y=�6��\v�N��dn(�:��6k���4^e�de�OxT��W%�����&��gs���֟+D;�&ӆB�G��L�i�<'��3Pͧï����މهP�%C��oS�f#*��I�!"�!��].�UM�$��W�7��s.�)$��+O������Z�Q]6�H5<�(H�L���w�l�=�@����-c=s^87��0�$��F{1�zYZ�B�@�3���N��0B�7���=\�8���a��i����(dʂ�qw����W5�+k�;ɊIݣ�mݽ�� ��!@�����%�8�A) �!7=��<5��.��Ӡ]ƄX���9AY0+= Μ�/k�-�}+�����F�"I$�B������荛��P������{��Z�֭��V�6u[,�*ʽ��c&o�Y�D>^�f<�X����:f�n��*]�b�ldo���.���c�
��ܜ|��{���<rd�D�Ȳy�Q9oU�<��/o��d��y�����W��N&o�Z=yX��s"q��0�&!!%$� C�O��6��i�ꚜ\g�*�]�|�#��'�)���Cy��Q�U";W����s0Z����QA���9�f^��2�N1�$.�T"��2P�#�v�tb�$1LH���+��yյ�����M�`��)-`�!4�5<��B�'vߴ ̖Ro�+4_kj�	��Z�ER�ٗpX)5˸�/4�x� 딒L�п{s�&�hA��.}��%�Kf����Ӭsݍh��K�%+�B���S��	*Ba����{v�k���ǠD����#k�X;̶+��LJS��|���]������b��3Ij�]�cJ�Z�Zg�ܝ{��͍w�]�ު�C\�מ�� �|U%[AZ���M���|xX�U� a�V��7I�qU��tK���иx�N\�L����3Dάz�A�~���?���ς�&#A@�(��E!B�J����<x������'Ql�w�T
��Jt+�&j�cd�O�]߽�%�u�ܷ>tL;��B�#{C�y���Y�^�o�Y�E�{dfb#�=�-�2��e��Ȁy<2P[�����QP�A�)���tJ�����r*��۾��D=�����y��I$�!'�s#��?�&.�vg2��!��|�!/#�"����Ș��l{!]�ǵ
��dKI���I�QyQ"��v(D���{�ꉍ��n�Pl[��C־�Lk���Thx��u��H�0��$D�
0A��u��ֺ�����9֔ZѽE{m�Xvyd�ɗ��G�^�t���AQQ)Q�dm���w�$9$r8�G�fv��g��z���܅�U���kUԸ��u�2G�m�`bq��j"E�DDbL1��E�m&fQD�l����/=�ëW�P�U��ʯ=m�L���#m�9��L�9���F����#Xg:�Ύ��^b<�S�ti���
3C�,w1P���ܹ��y����yK��έ���=�fUh��Y��0A޴m�ed�s�9�pT`�3u�tjg�7@wG�33&x�tD�>������Ӄ숹�� �>no8ۯ\��aU=7$�e�y�����><�cQ�=r��ȍ>D=��u�ǽݑM��hzdKZ �kx�D��r�-7�7ޞ9�HL(��I$�W��	�q�1�2��������u����w����at`�B9	�6!�<���m+�m�b����7��Csa
�'z7o&��uds62DA���!([{�E�{�A��3�ސ�dfl,�׺��3!l�·�;8�����JO�$q?��(��(����D>_�4s��	��u��M1� ��?�>���=#��8Y��x�M�y�;އSc����~�d\kU�`>����f�!���H���DI(�_v�t�2��S*���i���u����Ȗ{��7"{���ov���w��Һ�ϓsO��;��-0����b���<���`x�UN0Q���BdL��A�H[�{��z�nc�8���`��D#��r��Tr/��A(�%b���iN_Fy'jl��тQ(-�p��% 6�b�{^�D�j�����J�~PB�c��j.�d�L]����5�� ���nU��j�6G���0��S�V�� ���ERJ�0��S���ݧ�A�b ha!�~���|�|��u�-<��n؉��C9�l�F3#�=��B�h`��B)�%"J�"�����!�Ss�a�~�<�cO@Y�w���5�>݈�Q�8��F�#X[nL�0���5���êZ�H���@��`,7�_n��=�~{�� �"X�9 օ��qЄs�q
=�{����ׂeo���<JL��&1�3�ko[t�A1�����WZյ3��l�֤�.J���-,MξE}l�*���(-~��BuY�t$�0��IIFg+9]�Y_bj�W�P�XKyZ����{hfT7��Pu\R"N�<�I����ȠW{{�.�ڼ������K�w*�z2��O�sw��za\�~����J�m�9�L�����9�~������p�8��vL���8��?��~��t��r�� �2�Q�(����0�<��"d�O�W�]ͅ_c�ik�t��z���١&���@���Uy���z�誶��P�� ˮ��G���"�vJ���7ޏz��!.�I$�lJdU=Y�e�V��y��Ss�~cog��U5���9>'���A��C�8�~�����ަ�Oh�ׅH���<��u��m���E�e�M՗y�{��!Si�vy�?Â�<�I�ߵoK��-�b6��4��h*v��sgg8ɛ�6�WW�5,�A� ���'j�l���t����6]~����1�B�[����?�����-[0�8�0�qh��p�������~ə�9�s����Zc�tdG�}���𧧆��H��B�l��1
������kIb�uo 9}��y�Rۧ��(D#�
�����]�]x���ev˦�T�m�by���B�r�/�AQy��Ty
�G(�q� ��ƞ���h�cXCS�L�h��~�]�:�6��؁N��k@;<9�1�0�R�~ة�e�lO]����iP.z��ð�]��4�窨d7�r�jYh��8�#7����aJ�R[�veӫS�W��
|���B�Hj�zk��#�c���*�e��T����=\���ETE��,-LhӲ�#@fucWl�"�ɪ1jGV�{<�y{�2��(��[Z����cJ�������W'r,{�F�������8W�"ө�,�h:TF
�]$c"���ڴW�J���;nm�DZ6�m��m�6.(�E���^�5���,��B��9P�h����;h�uB�F��$m����d�6j=��[�*�����9:�{�֜,U���#��h����UF�y����ӊNMm��D[Q����l���ӵE�jF
�@�4�SD�-�;mwd�荋��bp�Ģ+��93�/r�yN�q��0��r%A�ՕɁ��J�r�*�U��[jȪ1UUQ���TAmUUTD���l������]E�Τ덗cX��҂��d�^��9����GLQ�iUz���yꪣ*6����*8W�V�G��v�sշ�m�5KO��y�)��f�p���h��<��PDF+��y�������tb�.)�Y�2	��{���l{���۸���ڕƌ�V�)sf^���'vr!j�bmK��ܧ-�Z���LbM�0�>�Af���Ѧ��Ӆ�\j�ȸm�R��k6�ɇ��(����1�/n��ȈZ&��'Lٸ�7p�;��C1C������ݿN�����7�ϘX�Y�4�qS��'y��8�N��dݭľQ�d�����j\5��fV�m˕�.Ys�K<�c�����<�)��{}⮇�{���ej�7y{{g��2���jq�2��[�isfoo4��U��اm�]��Ȼ��&�f�ԍ���������a�)��	K˼����x�{�R��BH���b#��M������r�DG���3���9�����u`��ѼYa-��/,G�.�3ɻ:ڶۍ��j �F�d�S����^.�FuCDD[Eso1C��)]PTU�v.Q�0z��Q�UNjT^�TF��V����""+�iX���j&B�&3[im���-�j��cGV���:��k�<�jDF-V���Vp���+�*��u��/�*�[���r-�"���rM��DEV1�9�[&����/U{�9+�ڌ��e�DDc��5DWm���.�[c�04,����Pʹ����ɨ�#j+�[l�gW�I��'`�N�+j�W����D�""!��DE-Q㻖�8W��U�vUs�e�P��.\=S@b�w+�V箊��^�um��v�ڈ�X��;[s9y�^ȥuDDH�DD�KN�S�?�VF��"�����Q�syx^�"<T�a�8V�F��toQ��r�eS�Ԕy{�U^t�6���w7w#lDIr.�h�����+ʪ	�R�b[m�FA$�2xff�����L�?��F�٦�"�����mf)^b�u�7nj�f���VQ�م����̊���Ƭ�����˜�Fd���Go�b�f�,�k(vc�}ϼ���c4���!^�����0�>f�CI�*�,�ٛo���&����A����/~&��s�y9}+�FTkm�7ym-�����4��r��p���.2�,���[Y����o�.��X��YF���e�4�J��&���<^�I��u�4x�����=x��[S2��`��/�c�-;������u_UV"���ݬ���r�Zr!W΁��-��Ŝ�P��{ўsm������wa��g��\
ح�ؿA}�@�f�{ 
�7�Z�P�@5��_E.	q&j9�SP糛Y�G O��=��<��B�B�@A0�L"h��-lub�	5��H�#h�X�3���93�<�h��vN^xE���rq�+E���v�es���<�<���-�����w{��N�F2�D�-p�&a2`S�t�<GUs����{*�$Q���
1��J�aܣ^TX���̱�9�N1ܵz'vM1�m��5��5k���7��U�U�)�pqX��v[���;���\���r!�su�ƭF���w��׶ՓM�ͩ}�Xk�Xe!)��5��0�'�;���wls���i�q���j�����G�� �����>����O�����D�,!�w.��צ�:X�VPޫ��A�A��A ��>.��{8�x%����s��B*�3��!h��˭���V��%s�B@؇����j��+����~�6���l�+R"�s���!v�q�E��]@��^�M��\�%i�mQ�z�Ǘ�v�rn���}�jZ��Ғq@��t�I)"�M�蒃�ް��V��n�\J'���|d<�e���ߩ>��� �B9����1�럶t����q�gp�g39:c��$�_����>Lx��8�!�L�z5P�;��=�8��
(����ʵ�ć�=5d��p1à���@�|��{�<�l�����c2�e�w�͵qz�p��9�Wƍ��e/���.��#�"��׼-�s�4�4����%��3������]d<߹x<z�I�QP�,�H��GC:�c��Ȫ}T@{C������qȗ�:%:-�3Z�@|Q����!����E��!��+����\N!ht6�����05jЛvO:��q4��^�<�=q]g#%�㖐G��`���0N�!�x��gd�w�</_B����(R汿צo��}�b�%�}>M��" �O���o�bE��E ���-�Í���ρ��丧�Br��W!����Z��6�O6��]Ӫ=��q��"ö��8�  �\A�6횽����&]��E����VDM��"��L�Bޭ�����x��:n�RKMH.II=BQ
(
��w�[���s�U�TL��u�K<��+�mt�g\�qm��D��F�T��~x�Wa��U{�g%����ּla�
�.��!�q�)���=�@�R'���	2_��`�� t�V���:bW�F� b$��2��F+]�`��.e��d<��ȍȆ7�R�@t:5�K���cU�|�垆x�u��s��m�$����"?y�n-���BO�Q@�(�Q �e{(p��3�N�s�s�	��4�&de=���a��8�@�(��}D7���&K=�p;��z�8�����R�a���7Z���LGs�9�;�9�J�j�U�Od��3a�!҅�ϵ72I�$Iq��˗�m�{�8%�@Ā��U�*o�D���W�Pօ��w��K~�V_D�=�W���0��;�Z���~����3q��A�R�
���8E k��������쩇�k��!e��JH�����sm5v��Y"��]Ǎ.z��f��}���m�r	��[���2Ys!���"�������cL�H�T��f��9��B���}{8��隱%�з���=��??��� �&�0�gC���X�Di���ɜ��p�d�p�'�_ߝ5�GK�2���wf!:��č.�[�����<�g���_���������.9��ȔE�ܚ�+��{��D�Y]=8������x��;-\NB!�r�AD*
�B0Z�2[��K��Vg�b��v7�G*\)�hyH�a�:V^����$�eU|�?Y��Sy {=b����Қ�2Pq����������Hy�`�N98�A�$<"o��(�x��W/<o�k�s�B"����5L��~ء���|"���	��� ��FNA�J�Kx@��"�gT`�Z��N�8s��&ts��a2�<�=c�*r��d�D[���M�@E#�ϟ�Dq��8'/���κ���T����)���]p����Hrb��>#A��ѴD���umS\��L;�cA��=��9�s����L�/'X�h���<9�ӌ<�<c�k2'l�#C=����9���$r��I E�;��
xb�o�V�*�w�u����\�]sc6V[oos����`eUX�y7g�gA�Ԭ@�kt4k��9�r�ծ\b�48DH��{,E,KA�b�� G�[�!k�A�6>�r�(�wz3Ӟ�lq3��{�9�A		0v�$?�-��x��y�}��m�r�1�+D�C^�@�)��//��~�k������Ҁ� �AIK`:�&�h�D�_���o�|�6������22��hlB@萑"'��k��N��R��*Z���ϺR��
��{���[��'uP�A�x�� $�E=Y�{��	��KIb���>�z%gdH�6ze^y�q}�d�|�����9�k�������!?	�<�4�b4�QE�'4�:h"f'����|>�p����_�F�(E�m�b���B)�'odZ�Mo�9���BDɩ���HH*GAռV[N!*�U�}���z]��hV!n��$�)j�0�8���d�Rz�痷�m^Uۢ�^�1����W׊%mn���;}1��t�]Sm��j�������ڗ���B8�d��h&�̘�.=�a.���:���צ`�����CQ�1��u���0�r��y����uw���{�DhU��D �������ݨ�w?^��(wOx�jy<�D
�~TAק�U۰d�tU6ڬ�!����9W"<�0��/W<�|(�I
Wfs��s�ՃA���;��WGs��u{�rpc�M�~_O�ϛ1 ������6�~�I�N�jK���=s7S����T�C��Ȱ�U��Ĥ�s�	XD��ݘӗ#L�O{i}�C�rU�zJ�=B��.r9��v�z��5
���Ă�P�I2�p��r$��}��M���8Ϟ��_^�B⸹"�6U������R�lC���[�b����.�6�n`��.�$�ŭ�Ei��b�fg��v��EP��n����|9�PPT ��rP]T+���.�zٟ��~��HB�o(y{�.v�z��n�\��z�TF^A�* ������k�����y�w�Ӣt�\��cە \��� XeU�`��H4:�g9�5L �d������B(��#(���,@���9���m�0ag}�=���6�T�K��{W)�#�+ѕ+�\J0ǱB*�<�18���!5�5�����՟e��O4�x5a��r"2P�[�I23^����A��A�(��&x��E��Awc�����}�xL�]�h���eU��Ǉts��(������aU�3�{�s����y &"R.�|������j�,����Sfꓹ��3��k����$��/Wm����C�l�xe����V=f�Ex�ܘ��y���$$a�G �P*e�3ț6����Ɵm��z�V�OJ�։[&��H����&??o����-��p�T�� `�| ���'���S�.Q1Z9�L�&Jf�4Dx��~|��|�B$@�B9�7hˢi�wiʰ���ĕ�6���Ώ2{�/��y����`�9�<��f{��H|�m���x��X
�Z"A/���;�p^����u!'��s�$Ր��_! ���6�9�/u�Wz:{i
��ᴡ�,S��xa�����݇��k׭Y$�s�v蔷Bm�ȍ�׫�ov������,Ll�R��"-D}�ǧ�SV>������Y{���:�D��#\=
�7LO�#���P���0`�� 6B���Ů�#K\9ףX�٭o��erǔ9NyW�b��eU�����X4�S�8y���p�r-��F���3ǐ\����I7�C
�S�.w�Җ���猐��O�� �}�'	Fb�8A5��n�rT펳/f��F�9�C9z��X���^Ng<`3
-墽�.y���s���m�S��t^���kJ�s�9�p=y!�s�]��^Vs�[3�G�Ljgf�s	�L��gkj�3e��2�6�\��U�m^�	�G�`�	> E�辉3�{�������	���D��6s���#߿�����3��A!��W��:��2*!S1/H!��i4����=���3S��%�@�@��r����Ը�����l��Q��Ҍ�D|UD�ɫ9��Ed��-<8�3	/���7`Ao&��U���
͗׵v�.�/�Q;Ӿ4[�$��I%$�!P*=-�ތ�W�EƱ�����D������ݔ�y�q��m��ǁ��̂ ��:'����yu���븯'��TOkf�,�,�����,���b qZÁ0�S	?�����a��s�d�գ��,��Ϟ���%�21C� �!�3\3՝W,�&�#ĺ�Ҵ�1�3냈��C{�jt �" �`L�P�lR��7��_�2�:t�ֿ� h���;3{��bհ�9���5��l�^֭ɑ�\2���護��g��\����{�����3=��:�o�t��:�G�v[�Bd�����q�4�{���nm�7@�r"+���+ݯ۠u8z`��{^���w��T�6\M�S�ҍ��z��v��	b%���uu��<����Ū�:�j����q� ��Q��"$���ݖhz{hڇ�^��$���ަ������b�� ��D>0A!�'edZZ�L@Ҋ袁@P�#33?�(���F�P���
�)�i�9o$���;���X���qN���ƅ�BA�;$�Bo�g�:z��o2�D��C1��|�:���C�Lə�^oL�E懳t����M!$m�A�o�h�.ؗ54jC���^�K*�4[��GՃa�+3a{�Sϳ�����o(̗b�\�i��]jmʱZv�wZ�ʼ�SqJ|eW-MƔ�U�"	ɸ}cor�)R#vm�/eV�hk����ɚ�lZ�����ƌ��i=Oz���	dg<��	^�tճ6�U6-��mi.����8;3kl�O;z�������{�cd�֌���l����!j�}!&{��:�!��}� �*!n�uY[s)kf���oV7[l�R6s=�<ӳ���{�ܛ܂�7vbaZ���D�6..�WV3d�/���:<䏭3-&�nkԵF>�뾬�=so�5�Tb�^K4�+<�J9���wgL�l<<�S�4hד��i�n���3s�7F�d�tj�fk�h��1iX��˛���k9���ފ>5�kث��dQ���{���}�{��D˓�ع��r����T��j�.ӨŨe�Vk9��q�U�K�F����71S��.��L�5SVϩl�W�j�W�-��<�5�I���,K�U6�<[k�ܶ�n[�6�����;���-)�Gۏ���k��b�����0<j:�b��Wnfv���+�!#@�x̚8�݋���Ƌ��ǭg��S_E/�6�w)��������� TD�I���R�$���MZ��9,�J���x�MYMX�KJ��Z��T��T�5K7WVcżL�#� ����W0@��r��|o�P��?L��Ȭ�%K�7u��î�ۮ<�,�Զ�.[W��g�C��������r	q��Y�Wv���c�%*'�Z�=�e�lm℺�E�<�ԙ���G�D�� �deVo�G��W���-�N�+f:�y��:�����8(��͜��Ƨ�"�Q8�F}�	��k����/ݕ�3��g��8s�1�	�~F��YD�A2:">�p�ȹMz�����Gy�f_�gJ�P;��9O�,������.��.f}~�����a�)ۧ hE�D�EE¿O�;���ZhJ��8���]�t�kgD�iX�-�����R��&=]�.{5�����G��$�eS�fz��
�۬T����&��j�R��z�z��*�h�5v�N��q�My�D4H�T�uJ�3�ɘ�=uxf��;Y�8�FN3k�ռ���o��T��A�jxC����?���p��u��GL���;��T��o�@��3�|q<� ��LV0\��rg0�с���ϴ���c\��&s�2fa�p&SY�0�{��IFKF�� �~b��"Hv�j�T���N:c�:s".�w=8��Y9ׁ��yN�[ �HIIЕ�|���w=�o=1hu�<�nz���s(�ZݿCT�7�9�f)$�J*TЛ��o!����C8�k��s����y��`"9O3��9���@q"Ds�{1��[���N?��������z��z=�a�6�AJ���%&`�r�Ji�Z$�m�.�D��TȉQ/}� ��O�B�xu��a02A1��U
:��8��dc���X�]Q�����u䣒��G��3�m��m��m��ʽ�,ċ�y���y���TH�#�ՍM��`m��s��N�+��p~���/�'���8�="G�>�����ǒm�z��}w�ue�snL?�Db��DD Рƹ��R��8��D;<9�frf��^N`�2�ʻ���	��\��rsp��8S�/�Z��d&��F�s���CA��xNz��QW������������vY����;p�zeL>D��MV���mY��<6�e���dn�̜�(�"�4�2�9�4��-��K��;�v��s��� S�A���=��|8�L�HJ�����Q4�
9��j	tH�A�9�3!�CSե�� b���e!D3���;��|mz5Dun��#���zDn�y�ַ٬�3J�zX���� ;;g�
Ԁ��&�V)n碷�9����B�Zx�Jq��*�[!��w���u���g� e���d���u-��U�fB�"d����	I	ҐA$�yP�'��7�0���z�mq�����\�	zW�d�:!��10���R�����⚢O����ޜw��s��3���d4�1�&o����4�|��D��2��/�~�IOaA�3��wюy����\�VE�F
�
x���RN7�ۗ�!����W�U�,�fU:�q"�k,��e��������o�f�x�O�\���.nN:���侹��cC�9�w`H��똴G*��C�9P�03�o�=�xÆF�D�&�z��o��eD�j�m������'��J��CWw�)G8����D�Bw��[����B�t=�
��	�xG��(�̅��l�c	C��A!KM~B�<�otۣ�s�\�~�D쬍@����w�B����TB(��2�B!è	�I���w�o���9̙�L8L�c��#��}��S���8Ar/f*�<�u�/ک��@m�����z���e�h-�;�i�N"�U���L�T���Bvﮢwf6�{�K(Z�Ut�J����;��bR�D�Ȑ�A*�KL��W���b��w������v�m���Z)�.�(��z�7���v�`yg�y����>��Z��\�Z�}�����Vj�|x�~�@,�2�_>��㧈HX
���w��=�5�v�	�T��[B6{c�	����J��9'���D}wm�Q� ��$�Bg@�mA��_7��˘X��`���	��BxB�u6��bh���rg	�94*1G����������7����fs��4�8������I	 �BBzz���q:��P��ũ<���<�-=��'>��>���9��w��#�q��K/��(��ш�6�����!�Mp�/��x���9�D	Aw�����g��S�����uC%�!�����ly���$�#��i�6V����.��uJ���*|&�!�8�9E���/^�O�ez�'+u�auw7jegW%�#����*Ep<�s���׆����C�;�V.P�kmjS���R�UO��ٗ}<~��\t|��L>0rA�B��&�{�cU�'x#[����D����+�M8a��"a���9�Φ�0c=o��{�>���9��u{C9ə�:t3-����!e��#�8�V�yJ��B�t�e�6�^E��!m���}��]N�5��)�w<9r:��C�βT5�����H:U��^�<;�*�WB�9���w�,(�]Ue-�4�~D/P��B�����zs��Pk�{\(7w.��4tJJ�&QA,*Y�ݏ��'zk����	bz��-�h"ڠ�m��=���N�����&I"ny{k��zM�Bq��o�bwG\����U,�޿R&^{�=CC��B�,Fa"h#� ���k"Z-�h3Q�"0k��tV���9�3�2�`zs��ZNy���6������'MTA�S �us��{4��s��t���K�4��e��f�V�{w)�%w*���/���im�YۛU�	�XH "��&k�5��ǰ��,�(���#���ʼ���i�;1E�x�S����l�xi�{�+�=&x�
Km%D[
���=�G"�<�Dy�0�r���<�EշO6V]F�R�󿨾9uH~��Km�Z�^<�E��+�\w�s#�QE�2Α�a	��w�{G&fs�DɇE�:Y8F:��U)��KGH
���@������Tķ�r�F)c#�.����b�zH4��I$���"S4��pH��9�Ѿں��gZ�oV7Y�� 2�4u"4y�Z�=��[RY�Ȩq)$��!*�������1�t6P �<s�����pNw��>��<��B���
K$���RHŔ2�z1��ڃ1<kY�jx{.1��-�T����b�׮D9t�0�8�I =�)5��<Ű����.՞�&��z�k�W��lY�O<,L9�C8��Ή�0F3����������s�{�s�8rS4�$:�H��A.
���#I#:&끥����)���}��,mm�\��v�q,����g$��-�@�C"=�u����?y���e�7|�.�׸�M��9M�M�ܴ���P��Y{�0v</I5Ӷ�ױ�3��e\�e���;�����&o�<���HG��N	�c�g3�	�7�׷X���
2a�Ad��!4���d�yC�
�	܊�df�T�\���(���A��I.�Hn�p���=u~����
��j:ЯXN��)]�}�`Ol��j1�!�A��kl�A��T=�����s5s�y��Q3 o[m� c��6:rpD,#B1"�)� �Au�{�	���E��(�8s�S����<bt:"d���U�H��A�:#�;�ȇq���=a�҇U3M�41�f���qhl� �[��P��G�hm�>�DC4���l����l�Ҝ��R5����b�_��4�o�2�FF�"1�CUy�TdCٔ�t�{�7λ�9U���]��nY��x\�`��9a��%︮|ͥm��و���v]�f�|ɝŝm6�v���me����։Z�\W��/&�:#�9 ��K+�3u��۞pOLyԎA�!��"p����ѹ�א(O���S*�(��=$kH`�mZ��NUBwD;�����z:�8����� ��}Hv{t]�ˑe���� tQ��`�Ho�0!>�;4a����QE�ES&M�c�8c��|8�g�>�����h-���p@n����o{g;ˁ�^��8�A$D@B@�]-·j4���r���ˋ7�'�{�^ C�� ��گ��o�o!8`r?�!H�Q�t{��P��.�������.{��bz���/�k��B��Y�<�JO�9�H��;��z;�e���;���� ���p�K�ٛ��{���z^��KE+��̾��Oؒ��<�
a/��.UB��R�b��d�p�������^4f�O�����U�?y����s�	.A�l���f�=���͐��P�Dn�����4o�����9��	�&���������}�w���0�����L��A����x�}��O�#��D�ԉ���hK�s��Si�}�l���h��r�a���I!$��%U	}�A�nǇ�TÛ��(�=��V�DD�2���{�b��y��p�b� �X��}�9�b�n	���
������kOXW��|�/8WV<�8pK�x�H-P5�.�̪�������k�~
q�F�Z��d�t��=�O_�c�%��`\,���"K<$���LGMGC�{:�<�s����9����a�_��!���)�C�eb|.n&W*��UUU��l�͘l�t�>g�f���x�QL��tT�f���~�И�)��,,.��m�.P��A���%��]Š�Pm��cu2�l�6�ٶ�f5f0��Ú�
��S0Z6�[m���+f̴D@�1E�"(����b*�(��*)��*}.psT6���<�dQDm��,b��TTi�,b���+��LEcR�"#LA�`�6L���S6ڠ	lAD$U�EP)b-��U )`���`��-�E!T���T4(��K�P<h*@'j`$;�@������R
TT1�PLT)@n�E,�P�D�4���P����ҊH(8�@K�TY�T&Ɨ#l�d�bCd��6�!��� �����ca�M�o/v@?�v����C:��M)��R�
�Ė����K?�@ B
lf�͆�V�٘kJ�614�F���%&���C?�)_o"�t�Ř�\�g�9��(��y��
�g�J�gB����W���~г8�G�t�B�������z�6j��e?Pu�x3���ߥI�EQ���m�H�
����?@��vk��Xeq���@�-�k�=�)v�6�����>���\o�f3��z�|"�l��~9,I&��R�� ������s���ì8������	��?���⼀<��U�q���e������O������?>�9Ǜ�6m��}�?G+f��?�������������׫x�{�����������iL!#��%��`O�L���y9�n�ﱟG���#��&���7���q�����?��.{7�[MI�OHTv@PY"cll?��*�@����<@e?~�}!���>(��!`�@j)�F�&cQ�")��m�kf6P�%ԤDA_�Q8�7Pي��v�oلyf�����3�65�93m�A���e�ٱ"�H"�H�"��ɖ���F$��4��[�M?1R��^e���
��6z�NB�b�K��[г37�Co8�dղ-L ��#��B���?���P����hZ�	���D��D���/�U"i���m�	�AL��_S!rj`p�
��q�TY�0�=Hs����	�����O�����7���kL�Mh��YH�A�Y$D�2"E�,�&�$I"Y&�K-4�E����%�%��M"E��H�k$I����Z�d�i���&��E�i�H�"KHK$I��i4�-�4��X�I�Z$��Yh��im,��Ye��M"Ye��md�id�K"�I��4k$B�-�I&�"�D$�&�k&�Z[HH�i�Ye�����i�Zk�$Z�L�-d�h�K$�Ĳ�H�H�Y"[D[Y,�&��bIe��$%��E��Z$�,�,�%���H��I�Z-�ɵ�ȖH�ki-4���k%��Y,�%��$%���K%�DD�����e���M$��D�M"�K$I��E��MH[[%�"�Kid�Y"M"�I��H�"%�b��"�K$�I��4�D�M,�Z�,L�Yd�E���kDX�D�M,���me�Mb$��Ye�����%��i��M-�-�d�Ie����d[Y6�I��I"�I�&�&�ie��ZYdYK%��mdE��Y%��dD�E���d���H�K$H�K%��i5�kh�K%�2E��D���Yk-��Zi�E��-�D��d�4���Z�-�DK-dE�d��%��e��M"�K%�kId�Y,���,��Bi$��dY"&�e��-��-"Ȳ"E���kH�I&�H�H��Kil�K"-dY,�֋DY$YdZi4�,�Yd�KE��2�[B�Yk$$�e�d"Ŧ�ZɢD��Y&"m,�I��M$�D�Z�",�K-d�$Z�ɬD�,�DK4��H�Y"D�Z�m2��,���"D�Yb��Y,��H�Zil�$$Zk�D�e��%�[Y��K$�I��%�%�$I�-&�k%�-4�d�ֈ�%�[h��X��dD�!$�,�Ke�E��m,�D��Mh�I���E��M2$HZ�d�E���!&�&�I��X�H�d�H�Є���d��m$Y,�"$���h[K!Z�4�K!d�i�%��"�H�d%�$���X����I�d,�ֲ�K%�Y"Œ%��,�E�,,�KbD�Yi"M"Y,�,�&D[Ik$�$I�H"�Ikh�Y	�M�d�e��&��$Kd�D�,����D�Y,��kY$&�XY,�B$Ym"�$X�idY&��iE�$BBD�,�-d��&�[%��d�d�e�Yk$�,�Z-dYk$�$I&���4�Y,��d�IdD,�KiYm�F�ID��,���,��Y,�I��"Mi��Y,�%������dE����d�"M"k"%�d��E�-4&�%��,K-d�M$H��K��[KkYh�K"�D��Zd�dMe��m,�D��Y&��im,�K"MY&�4H�-	4�I&��%�&�4�"YdKZ%��d��d��i4�imE��!h�hH�-%�ċY,��E��$�Z%����H��i�I-���!bɭ�K%�d�i5�-���D�[Z�I4�D5��D��		"-4�M5��K%�,��!,��YE�Yh�Z�D�K&��Zi%��,�,�H�I�Z$�&�$�%��H�$Ki%�K-YmŖH�-���&�&�YdI�K%��I4�Y,���4��&�Mh��f�,�Z��K"YmdBD�d�$K$��!m�-K"�d[H�Y4�$K!Y$��$���	$�",�Z$K-ȚD�Y&�I�K-d���-�[B�d�&�%��"�dE��%��4��Kh�D�me�K%�5��[i�B,�Yd�Yk#[Z$I��m,�K�E��bM"[Z�M"Ml�Y$�,�$$��"%���Ih�Z�5���d,��MdD�Yh�Zi5���$���E�%���"$�d��M4Z�[kD�"Diie�k$I��̑"H��Z�Yh�Z"�e�,�K,�h��"�e���I�Z&�Yk%�D���I��&�"�id�k-��i,��H�I$�e��d�Y&�H�ZK$�k[E�d�ȖZ�4�5��d��"ki�$�&�L�ֲD��e�mkE����K-4F�$M5�K%��D��5�m2BI,�Zi4�,�L��$�-e�D�k$Ki4��X�ZibD�d���ɥ��E��e�D����KIm"�Y$�$%��KdE��Mkd&��Z�Yd��D�-��Ye�DH�i�d�D�Y�"-��-e�X��$E��D�d��I��ȲɤI"&�2"�M"�H�I,�-���e�Z�4�YD�"MK$%�Mkid�%�i%�Yh�H�Z,���"[DH�ֲD��Y,��&�K$֛K-,�Y"[H�,�D�[Y$ȚZ-dY,��	I��$�il��dY"KD�"D���ɢM-i��e��H�K$ȴD��-m"E��Z�i��Y,�H����Z�D��e��&�K%�$�Iki��Zh��ֲ�i&̒�d��K,�M"h�I,�,�I��h�,�$���D%��e�Y,�kH�Z�e�	��L�Z$�kD�YMH�K�E�,��d�%��"�$�"&���D%�4��KKkB-�YdMh�Yf���$�D�Yh�k%�D�X�Y,�H�e���ȲI�%�$I�"�I��id�Ml��,�։%���kD�L�K$K-id�D�Y,�I����Y"���,�$�-���E��-���̒[m&�K1-��$�KlKa$�Ka&�F%�I����I�,ĒM`�!�m��֛,�"̑��m$[h��2[i6K2M�2�ͤ��bM�m�ؐH,�i�I,�,�Z���Z�ȲD�&�h��Ye��&�5����m��KD�Mdք�k$֚ɤ�Z�d�d�Y,�!m���dkkYk$�e�"M$��-����Y4H�,�ZI!"M,�HI���X���4�Zie��Ymk$��4K%��dY�$�HK%�$K%�$֚D�K-�"!k,�Z�"Ȳ�h"�dE���٭�̚ȓY%��e�K%��K%�Y5�d�KY4�X�,�&�,�Ie�ȵ���"ie�HI$�2�"Y"Y,Z�-�-5���M,�"M,�$�D���l�M,�,�M�Mk-����d�i�I���DYL�D��H[DY"Y,�"Mh���E��$-iD��[Zie��$I����I"�I�M#K%�M-�ɴ�!,�k-�Y&�I%�Z$H�D"-d�,��Y"[D�DYH�%�H���D%���HYd�ȉe�4��D�F���e�KidM,��I&�$�d�Yi�D�B$���e��I��d���-�&�H��h��[M%���[Y!"Yk-��D��X�m��I��%�I	�M,��-�i��X��H���,�Y"�"�$HZ�,�i�-�-����Yk$I��"kYdI&�!�D�lY,�$��d[Yd�"��,�Mm&��Z%���e��h�б$�,�,�M�5����D!h�I��"Y��I4�Y&�&�,�i$�Z�[Mm",�I���Ie���4�&K$Kh�%���-���4H����e�"�mh�Z�Y%����Y"D��E��%��,��Y,�k,��ɤֲMe�i��5�ZDY�"%�%��$K-$֋Mi��YhH�HX��k&�%����f�̑5�&Z$B�d�&Z$��d�D�k-d�Y,��H�2k&�I��e��3KM,��E���։e���BM"E�B$��I����D�Y,�-h��șd�D�"k-�ֶ��Zi,`B"A�����m���C �X�D}s�����MZ��� 5������Z��E?�{A��a����g�+_s�=��<��#�o���5�n~+�/�?b��:>���?���ӡ��
�(���F�1��0Cރ���2aݩIh�о�5xJ�|ƙ����;;U�  `��ב��҈*C��PP��O��0����O�j���8(?�a�Ћ�?P�_A��	�~��31��6y����Hs���?@r��
?"*�1�'���:<����hϴ�fޟ-��>�?��F���P��� 2��C9�~��*�[AA��4?��t6��5yR��?�~�?�c�d P��D?8B�!ʃ��	P�!�_��T��K����`8�����r�����~?����㕝
�"��_�mKr�jgi3���F���% 8-�$-��h��wi����SH%���M#�#�A�&H@�c�"��S����!��������X�G*�P��?��\���?�O��XV���*��?���(~?���@T@
�����\�/g�3�_��^��R�4��	H�0HU`"��Ѝy�GYuӉ�\n|��X@�+��)�!�(B%�0c���O�L ���D�������]r��ަ@,+��������K����c�2��d����rV���o�TEzQ��q�'�c����*�Ϗ��� ��_�+������wU��σ�OЂ=?���d!�~���� p�#����B��ʬ���GZ�7��01�o��yf=�>��ρfL�c~�ѹ�<�a�"�H\�<W��9/j�r�����~� �x�?�0?jE�W:q������sA���)_���$��kw9�=�H���ONS�3��
bbz�B�����?�C������]��BBob �